//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename:ipsxe_floating_point_log_32_axi_v1_0.v
// Function: p=ln(z)
//           zsize:z > 0
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ns

module ipsxe_floating_point_log_64_axi_v1_0 #(
    parameter FLOAT_EXP_WIDTH = 11,
    parameter FLOAT_FRAC_WIDTH = 53,
    parameter ITERATION_NUM = 3
)
(
    input i_clk, //aclk
    input i_aclken,
    input i_rst_n, //aresetn
    input [FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-1:0] i_data, //s_axis_a_tdata
    input i_valid, //s_axis_a_tvalid
    output [FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-1:0] o_ln_float, //m_axis_result_tdata
    output o_invalid_op,
    output o_overflow, 
    output o_underflow,
    output o_valid //m_axis_result_tvalid
);

//look up table 
wire [52:0] f1_rom [1023:0];
assign f1_rom[0] = 53'd4503599627370496;
assign f1_rom[1] = 52'd4499201580859392;
assign f1_rom[2] = 52'd4494803534348288;
assign f1_rom[3] = 52'd4490405487837184;
assign f1_rom[4] = 52'd4486007441326080;
assign f1_rom[5] = 52'd4481609394814976;
assign f1_rom[6] = 52'd4477211348303872;
assign f1_rom[7] = 52'd4472813301792768;
assign f1_rom[8] = 52'd4468415255281664;
assign f1_rom[9] = 52'd4464017208770560;
assign f1_rom[10] = 52'd4459619162259456;
assign f1_rom[11] = 52'd4455221115748352;
assign f1_rom[12] = 52'd4450823069237248;
assign f1_rom[13] = 52'd4446425022726144;
assign f1_rom[14] = 52'd4442026976215040;
assign f1_rom[15] = 52'd4437628929703936;
assign f1_rom[16] = 52'd4433230883192832;
assign f1_rom[17] = 52'd4428832836681728;
assign f1_rom[18] = 52'd4424434790170624;
assign f1_rom[19] = 52'd4420036743659520;
assign f1_rom[20] = 52'd4415638697148416;
assign f1_rom[21] = 52'd4411240650637312;
assign f1_rom[22] = 52'd4406842604126208;
assign f1_rom[23] = 52'd4406842604126208;
assign f1_rom[24] = 52'd4402444557615104;
assign f1_rom[25] = 52'd4398046511104000;
assign f1_rom[26] = 52'd4393648464592896;
assign f1_rom[27] = 52'd4389250418081792;
assign f1_rom[28] = 52'd4384852371570688;
assign f1_rom[29] = 52'd4380454325059584;
assign f1_rom[30] = 52'd4376056278548480;
assign f1_rom[31] = 52'd4371658232037376;
assign f1_rom[32] = 52'd4367260185526272;
assign f1_rom[33] = 52'd4362862139015168;
assign f1_rom[34] = 52'd4358464092504064;
assign f1_rom[35] = 52'd4354066045992960;
assign f1_rom[36] = 52'd4349667999481856;
assign f1_rom[37] = 52'd4345269952970752;
assign f1_rom[38] = 52'd4340871906459648;
assign f1_rom[39] = 52'd4336473859948544;
assign f1_rom[40] = 52'd4336473859948544;
assign f1_rom[41] = 52'd4332075813437440;
assign f1_rom[42] = 52'd4327677766926336;
assign f1_rom[43] = 52'd4323279720415232;
assign f1_rom[44] = 52'd4318881673904128;
assign f1_rom[45] = 52'd4314483627393024;
assign f1_rom[46] = 52'd4310085580881920;
assign f1_rom[47] = 52'd4305687534370816;
assign f1_rom[48] = 52'd4301289487859712;
assign f1_rom[49] = 52'd4296891441348608;
assign f1_rom[50] = 52'd4292493394837504;
assign f1_rom[51] = 52'd4288095348326400;
assign f1_rom[52] = 52'd4288095348326400;
assign f1_rom[53] = 52'd4283697301815296;
assign f1_rom[54] = 52'd4279299255304192;
assign f1_rom[55] = 52'd4274901208793088;
assign f1_rom[56] = 52'd4270503162281984;
assign f1_rom[57] = 52'd4266105115770880;
assign f1_rom[58] = 52'd4261707069259776;
assign f1_rom[59] = 52'd4257309022748672;
assign f1_rom[60] = 52'd4252910976237568;
assign f1_rom[61] = 52'd4248512929726464;
assign f1_rom[62] = 52'd4248512929726464;
assign f1_rom[63] = 52'd4244114883215360;
assign f1_rom[64] = 52'd4239716836704256;
assign f1_rom[65] = 52'd4235318790193152;
assign f1_rom[66] = 52'd4230920743682048;
assign f1_rom[67] = 52'd4226522697170944;
assign f1_rom[68] = 52'd4222124650659840;
assign f1_rom[69] = 52'd4217726604148736;
assign f1_rom[70] = 52'd4213328557637632;
assign f1_rom[71] = 52'd4213328557637632;
assign f1_rom[72] = 52'd4208930511126528;
assign f1_rom[73] = 52'd4204532464615424;
assign f1_rom[74] = 52'd4200134418104320;
assign f1_rom[75] = 52'd4195736371593216;
assign f1_rom[76] = 52'd4191338325082112;
assign f1_rom[77] = 52'd4186940278571008;
assign f1_rom[78] = 52'd4186940278571008;
assign f1_rom[79] = 52'd4182542232059904;
assign f1_rom[80] = 52'd4178144185548800;
assign f1_rom[81] = 52'd4173746139037696;
assign f1_rom[82] = 52'd4169348092526592;
assign f1_rom[83] = 52'd4164950046015488;
assign f1_rom[84] = 52'd4160551999504384;
assign f1_rom[85] = 52'd4160551999504384;
assign f1_rom[86] = 52'd4156153952993280;
assign f1_rom[87] = 52'd4151755906482176;
assign f1_rom[88] = 52'd4147357859971072;
assign f1_rom[89] = 52'd4142959813459968;
assign f1_rom[90] = 52'd4138561766948864;
assign f1_rom[91] = 52'd4134163720437760;
assign f1_rom[92] = 52'd4134163720437760;
assign f1_rom[93] = 52'd4129765673926656;
assign f1_rom[94] = 52'd4125367627415552;
assign f1_rom[95] = 52'd4120969580904448;
assign f1_rom[96] = 52'd4116571534393344;
assign f1_rom[97] = 52'd4112173487882240;
assign f1_rom[98] = 52'd4112173487882240;
assign f1_rom[99] = 52'd4107775441371136;
assign f1_rom[100] = 52'd4103377394860032;
assign f1_rom[101] = 52'd4098979348348928;
assign f1_rom[102] = 52'd4094581301837824;
assign f1_rom[103] = 52'd4090183255326720;
assign f1_rom[104] = 52'd4090183255326720;
assign f1_rom[105] = 52'd4085785208815616;
assign f1_rom[106] = 52'd4081387162304512;
assign f1_rom[107] = 52'd4076989115793408;
assign f1_rom[108] = 52'd4072591069282304;
assign f1_rom[109] = 52'd4068193022771200;
assign f1_rom[110] = 52'd4068193022771200;
assign f1_rom[111] = 52'd4063794976260096;
assign f1_rom[112] = 52'd4059396929748992;
assign f1_rom[113] = 52'd4054998883237888;
assign f1_rom[114] = 52'd4050600836726784;
assign f1_rom[115] = 52'd4050600836726784;
assign f1_rom[116] = 52'd4046202790215680;
assign f1_rom[117] = 52'd4041804743704576;
assign f1_rom[118] = 52'd4037406697193472;
assign f1_rom[119] = 52'd4033008650682368;
assign f1_rom[120] = 52'd4033008650682368;
assign f1_rom[121] = 52'd4028610604171264;
assign f1_rom[122] = 52'd4024212557660160;
assign f1_rom[123] = 52'd4019814511149056;
assign f1_rom[124] = 52'd4015416464637952;
assign f1_rom[125] = 52'd4015416464637952;
assign f1_rom[126] = 52'd4011018418126848;
assign f1_rom[127] = 52'd4006620371615744;
assign f1_rom[128] = 52'd4002222325104640;
assign f1_rom[129] = 52'd3997824278593536;
assign f1_rom[130] = 52'd3997824278593536;
assign f1_rom[131] = 52'd3993426232082432;
assign f1_rom[132] = 52'd3989028185571328;
assign f1_rom[133] = 52'd3984630139060224;
assign f1_rom[134] = 52'd3984630139060224;
assign f1_rom[135] = 52'd3980232092549120;
assign f1_rom[136] = 52'd3975834046038016;
assign f1_rom[137] = 52'd3971435999526912;
assign f1_rom[138] = 52'd3967037953015808;
assign f1_rom[139] = 52'd3967037953015808;
assign f1_rom[140] = 52'd3962639906504704;
assign f1_rom[141] = 52'd3958241859993600;
assign f1_rom[142] = 52'd3953843813482496;
assign f1_rom[143] = 52'd3953843813482496;
assign f1_rom[144] = 52'd3949445766971392;
assign f1_rom[145] = 52'd3945047720460288;
assign f1_rom[146] = 52'd3940649673949184;
assign f1_rom[147] = 52'd3936251627438080;
assign f1_rom[148] = 52'd3936251627438080;
assign f1_rom[149] = 52'd3931853580926976;
assign f1_rom[150] = 52'd3927455534415872;
assign f1_rom[151] = 52'd3923057487904768;
assign f1_rom[152] = 52'd3923057487904768;
assign f1_rom[153] = 52'd3918659441393664;
assign f1_rom[154] = 52'd3914261394882560;
assign f1_rom[155] = 52'd3909863348371456;
assign f1_rom[156] = 52'd3909863348371456;
assign f1_rom[157] = 52'd3905465301860352;
assign f1_rom[158] = 52'd3901067255349248;
assign f1_rom[159] = 52'd3896669208838144;
assign f1_rom[160] = 52'd3896669208838144;
assign f1_rom[161] = 52'd3892271162327040;
assign f1_rom[162] = 52'd3887873115815936;
assign f1_rom[163] = 52'd3883475069304832;
assign f1_rom[164] = 52'd3883475069304832;
assign f1_rom[165] = 52'd3879077022793728;
assign f1_rom[166] = 52'd3874678976282624;
assign f1_rom[167] = 52'd3870280929771520;
assign f1_rom[168] = 52'd3870280929771520;
assign f1_rom[169] = 52'd3865882883260416;
assign f1_rom[170] = 52'd3861484836749312;
assign f1_rom[171] = 52'd3857086790238208;
assign f1_rom[172] = 52'd3857086790238208;
assign f1_rom[173] = 52'd3852688743727104;
assign f1_rom[174] = 52'd3848290697216000;
assign f1_rom[175] = 52'd3848290697216000;
assign f1_rom[176] = 52'd3843892650704896;
assign f1_rom[177] = 52'd3839494604193792;
assign f1_rom[178] = 52'd3835096557682688;
assign f1_rom[179] = 52'd3835096557682688;
assign f1_rom[180] = 52'd3830698511171584;
assign f1_rom[181] = 52'd3826300464660480;
assign f1_rom[182] = 52'd3821902418149376;
assign f1_rom[183] = 52'd3821902418149376;
assign f1_rom[184] = 52'd3817504371638272;
assign f1_rom[185] = 52'd3813106325127168;
assign f1_rom[186] = 52'd3813106325127168;
assign f1_rom[187] = 52'd3808708278616064;
assign f1_rom[188] = 52'd3804310232104960;
assign f1_rom[189] = 52'd3799912185593856;
assign f1_rom[190] = 52'd3799912185593856;
assign f1_rom[191] = 52'd3795514139082752;
assign f1_rom[192] = 52'd3791116092571648;
assign f1_rom[193] = 52'd3791116092571648;
assign f1_rom[194] = 52'd3786718046060544;
assign f1_rom[195] = 52'd3782319999549440;
assign f1_rom[196] = 52'd3777921953038336;
assign f1_rom[197] = 52'd3777921953038336;
assign f1_rom[198] = 52'd3773523906527232;
assign f1_rom[199] = 52'd3769125860016128;
assign f1_rom[200] = 52'd3769125860016128;
assign f1_rom[201] = 52'd3764727813505024;
assign f1_rom[202] = 52'd3760329766993920;
assign f1_rom[203] = 52'd3760329766993920;
assign f1_rom[204] = 52'd3755931720482816;
assign f1_rom[205] = 52'd3751533673971712;
assign f1_rom[206] = 52'd3751533673971712;
assign f1_rom[207] = 52'd3747135627460608;
assign f1_rom[208] = 52'd3742737580949504;
assign f1_rom[209] = 52'd3738339534438400;
assign f1_rom[210] = 52'd3738339534438400;
assign f1_rom[211] = 52'd3733941487927296;
assign f1_rom[212] = 52'd3729543441416192;
assign f1_rom[213] = 52'd3729543441416192;
assign f1_rom[214] = 52'd3725145394905088;
assign f1_rom[215] = 52'd3720747348393984;
assign f1_rom[216] = 52'd3720747348393984;
assign f1_rom[217] = 52'd3716349301882880;
assign f1_rom[218] = 52'd3711951255371776;
assign f1_rom[219] = 52'd3711951255371776;
assign f1_rom[220] = 52'd3707553208860672;
assign f1_rom[221] = 52'd3703155162349568;
assign f1_rom[222] = 52'd3703155162349568;
assign f1_rom[223] = 52'd3698757115838464;
assign f1_rom[224] = 52'd3694359069327360;
assign f1_rom[225] = 52'd3694359069327360;
assign f1_rom[226] = 52'd3689961022816256;
assign f1_rom[227] = 52'd3685562976305152;
assign f1_rom[228] = 52'd3685562976305152;
assign f1_rom[229] = 52'd3681164929794048;
assign f1_rom[230] = 52'd3676766883282944;
assign f1_rom[231] = 52'd3676766883282944;
assign f1_rom[232] = 52'd3672368836771840;
assign f1_rom[233] = 52'd3667970790260736;
assign f1_rom[234] = 52'd3667970790260736;
assign f1_rom[235] = 52'd3663572743749632;
assign f1_rom[236] = 52'd3659174697238528;
assign f1_rom[237] = 52'd3659174697238528;
assign f1_rom[238] = 52'd3654776650727424;
assign f1_rom[239] = 52'd3650378604216320;
assign f1_rom[240] = 52'd3650378604216320;
assign f1_rom[241] = 52'd3645980557705216;
assign f1_rom[242] = 52'd3641582511194112;
assign f1_rom[243] = 52'd3641582511194112;
assign f1_rom[244] = 52'd3637184464683008;
assign f1_rom[245] = 52'd3632786418171904;
assign f1_rom[246] = 52'd3632786418171904;
assign f1_rom[247] = 52'd3628388371660800;
assign f1_rom[248] = 52'd3623990325149696;
assign f1_rom[249] = 52'd3623990325149696;
assign f1_rom[250] = 52'd3619592278638592;
assign f1_rom[251] = 52'd3615194232127488;
assign f1_rom[252] = 52'd3615194232127488;
assign f1_rom[253] = 52'd3610796185616384;
assign f1_rom[254] = 52'd3606398139105280;
assign f1_rom[255] = 52'd3606398139105280;
assign f1_rom[256] = 52'd3602000092594176;
assign f1_rom[257] = 52'd3602000092594176;
assign f1_rom[258] = 52'd3597602046083072;
assign f1_rom[259] = 52'd3593203999571968;
assign f1_rom[260] = 52'd3593203999571968;
assign f1_rom[261] = 52'd3588805953060864;
assign f1_rom[262] = 52'd3584407906549760;
assign f1_rom[263] = 52'd3584407906549760;
assign f1_rom[264] = 52'd3580009860038656;
assign f1_rom[265] = 52'd3575611813527552;
assign f1_rom[266] = 52'd3575611813527552;
assign f1_rom[267] = 52'd3571213767016448;
assign f1_rom[268] = 52'd3571213767016448;
assign f1_rom[269] = 52'd3566815720505344;
assign f1_rom[270] = 52'd3562417673994240;
assign f1_rom[271] = 52'd3562417673994240;
assign f1_rom[272] = 52'd3558019627483136;
assign f1_rom[273] = 52'd3553621580972032;
assign f1_rom[274] = 52'd3553621580972032;
assign f1_rom[275] = 52'd3549223534460928;
assign f1_rom[276] = 52'd3549223534460928;
assign f1_rom[277] = 52'd3544825487949824;
assign f1_rom[278] = 52'd3540427441438720;
assign f1_rom[279] = 52'd3540427441438720;
assign f1_rom[280] = 52'd3536029394927616;
assign f1_rom[281] = 52'd3536029394927616;
assign f1_rom[282] = 52'd3531631348416512;
assign f1_rom[283] = 52'd3527233301905408;
assign f1_rom[284] = 52'd3527233301905408;
assign f1_rom[285] = 52'd3522835255394304;
assign f1_rom[286] = 52'd3518437208883200;
assign f1_rom[287] = 52'd3518437208883200;
assign f1_rom[288] = 52'd3514039162372096;
assign f1_rom[289] = 52'd3514039162372096;
assign f1_rom[290] = 52'd3509641115860992;
assign f1_rom[291] = 52'd3505243069349888;
assign f1_rom[292] = 52'd3505243069349888;
assign f1_rom[293] = 52'd3500845022838784;
assign f1_rom[294] = 52'd3500845022838784;
assign f1_rom[295] = 52'd3496446976327680;
assign f1_rom[296] = 52'd3492048929816576;
assign f1_rom[297] = 52'd3492048929816576;
assign f1_rom[298] = 52'd3487650883305472;
assign f1_rom[299] = 52'd3487650883305472;
assign f1_rom[300] = 52'd3483252836794368;
assign f1_rom[301] = 52'd3478854790283264;
assign f1_rom[302] = 52'd3478854790283264;
assign f1_rom[303] = 52'd3474456743772160;
assign f1_rom[304] = 52'd3474456743772160;
assign f1_rom[305] = 52'd3470058697261056;
assign f1_rom[306] = 52'd3465660650749952;
assign f1_rom[307] = 52'd3465660650749952;
assign f1_rom[308] = 52'd3461262604238848;
assign f1_rom[309] = 52'd3461262604238848;
assign f1_rom[310] = 52'd3456864557727744;
assign f1_rom[311] = 52'd3452466511216640;
assign f1_rom[312] = 52'd3452466511216640;
assign f1_rom[313] = 52'd3448068464705536;
assign f1_rom[314] = 52'd3448068464705536;
assign f1_rom[315] = 52'd3443670418194432;
assign f1_rom[316] = 52'd3443670418194432;
assign f1_rom[317] = 52'd3439272371683328;
assign f1_rom[318] = 52'd3434874325172224;
assign f1_rom[319] = 52'd3434874325172224;
assign f1_rom[320] = 52'd3430476278661120;
assign f1_rom[321] = 52'd3430476278661120;
assign f1_rom[322] = 52'd3426078232150016;
assign f1_rom[323] = 52'd3421680185638912;
assign f1_rom[324] = 52'd3421680185638912;
assign f1_rom[325] = 52'd3417282139127808;
assign f1_rom[326] = 52'd3417282139127808;
assign f1_rom[327] = 52'd3412884092616704;
assign f1_rom[328] = 52'd3412884092616704;
assign f1_rom[329] = 52'd3408486046105600;
assign f1_rom[330] = 52'd3404087999594496;
assign f1_rom[331] = 52'd3404087999594496;
assign f1_rom[332] = 52'd3399689953083392;
assign f1_rom[333] = 52'd3399689953083392;
assign f1_rom[334] = 52'd3395291906572288;
assign f1_rom[335] = 52'd3395291906572288;
assign f1_rom[336] = 52'd3390893860061184;
assign f1_rom[337] = 52'd3386495813550080;
assign f1_rom[338] = 52'd3386495813550080;
assign f1_rom[339] = 52'd3382097767038976;
assign f1_rom[340] = 52'd3382097767038976;
assign f1_rom[341] = 52'd3377699720527872;
assign f1_rom[342] = 52'd3377699720527872;
assign f1_rom[343] = 52'd3373301674016768;
assign f1_rom[344] = 52'd3373301674016768;
assign f1_rom[345] = 52'd3368903627505664;
assign f1_rom[346] = 52'd3364505580994560;
assign f1_rom[347] = 52'd3364505580994560;
assign f1_rom[348] = 52'd3360107534483456;
assign f1_rom[349] = 52'd3360107534483456;
assign f1_rom[350] = 52'd3355709487972352;
assign f1_rom[351] = 52'd3355709487972352;
assign f1_rom[352] = 52'd3351311441461248;
assign f1_rom[353] = 52'd3346913394950144;
assign f1_rom[354] = 52'd3346913394950144;
assign f1_rom[355] = 52'd3342515348439040;
assign f1_rom[356] = 52'd3342515348439040;
assign f1_rom[357] = 52'd3338117301927936;
assign f1_rom[358] = 52'd3338117301927936;
assign f1_rom[359] = 52'd3333719255416832;
assign f1_rom[360] = 52'd3333719255416832;
assign f1_rom[361] = 52'd3329321208905728;
assign f1_rom[362] = 52'd3329321208905728;
assign f1_rom[363] = 52'd3324923162394624;
assign f1_rom[364] = 52'd3320525115883520;
assign f1_rom[365] = 52'd3320525115883520;
assign f1_rom[366] = 52'd3316127069372416;
assign f1_rom[367] = 52'd3316127069372416;
assign f1_rom[368] = 52'd3311729022861312;
assign f1_rom[369] = 52'd3311729022861312;
assign f1_rom[370] = 52'd3307330976350208;
assign f1_rom[371] = 52'd3307330976350208;
assign f1_rom[372] = 52'd3302932929839104;
assign f1_rom[373] = 52'd3302932929839104;
assign f1_rom[374] = 52'd3298534883328000;
assign f1_rom[375] = 52'd3298534883328000;
assign f1_rom[376] = 52'd3294136836816896;
assign f1_rom[377] = 52'd3289738790305792;
assign f1_rom[378] = 52'd3289738790305792;
assign f1_rom[379] = 52'd3285340743794688;
assign f1_rom[380] = 52'd3285340743794688;
assign f1_rom[381] = 52'd3280942697283584;
assign f1_rom[382] = 52'd3280942697283584;
assign f1_rom[383] = 52'd3276544650772480;
assign f1_rom[384] = 52'd3276544650772480;
assign f1_rom[385] = 52'd3272146604261376;
assign f1_rom[386] = 52'd3272146604261376;
assign f1_rom[387] = 52'd3267748557750272;
assign f1_rom[388] = 52'd3267748557750272;
assign f1_rom[389] = 52'd3263350511239168;
assign f1_rom[390] = 52'd3263350511239168;
assign f1_rom[391] = 52'd3258952464728064;
assign f1_rom[392] = 52'd3258952464728064;
assign f1_rom[393] = 52'd3254554418216960;
assign f1_rom[394] = 52'd3250156371705856;
assign f1_rom[395] = 52'd3250156371705856;
assign f1_rom[396] = 52'd3245758325194752;
assign f1_rom[397] = 52'd3245758325194752;
assign f1_rom[398] = 52'd3241360278683648;
assign f1_rom[399] = 52'd3241360278683648;
assign f1_rom[400] = 52'd3236962232172544;
assign f1_rom[401] = 52'd3236962232172544;
assign f1_rom[402] = 52'd3232564185661440;
assign f1_rom[403] = 52'd3232564185661440;
assign f1_rom[404] = 52'd3228166139150336;
assign f1_rom[405] = 52'd3228166139150336;
assign f1_rom[406] = 52'd3223768092639232;
assign f1_rom[407] = 52'd3223768092639232;
assign f1_rom[408] = 52'd3219370046128128;
assign f1_rom[409] = 52'd3219370046128128;
assign f1_rom[410] = 52'd3214971999617024;
assign f1_rom[411] = 52'd3214971999617024;
assign f1_rom[412] = 52'd3210573953105920;
assign f1_rom[413] = 52'd3210573953105920;
assign f1_rom[414] = 52'd3206175906594816;
assign f1_rom[415] = 52'd3206175906594816;
assign f1_rom[416] = 52'd3201777860083712;
assign f1_rom[417] = 52'd3201777860083712;
assign f1_rom[418] = 52'd3197379813572608;
assign f1_rom[419] = 52'd3197379813572608;
assign f1_rom[420] = 52'd3192981767061504;
assign f1_rom[421] = 52'd3192981767061504;
assign f1_rom[422] = 52'd3188583720550400;
assign f1_rom[423] = 52'd3188583720550400;
assign f1_rom[424] = 52'd3184185674039296;
assign f1_rom[425] = 52'd3184185674039296;
assign f1_rom[426] = 52'd3179787627528192;
assign f1_rom[427] = 52'd3179787627528192;
assign f1_rom[428] = 52'd3175389581017088;
assign f1_rom[429] = 52'd3175389581017088;
assign f1_rom[430] = 52'd3170991534505984;
assign f1_rom[431] = 52'd3170991534505984;
assign f1_rom[432] = 52'd3166593487994880;
assign f1_rom[433] = 52'd3166593487994880;
assign f1_rom[434] = 52'd3162195441483776;
assign f1_rom[435] = 52'd3162195441483776;
assign f1_rom[436] = 52'd3157797394972672;
assign f1_rom[437] = 52'd3157797394972672;
assign f1_rom[438] = 52'd3153399348461568;
assign f1_rom[439] = 52'd3153399348461568;
assign f1_rom[440] = 52'd3149001301950464;
assign f1_rom[441] = 52'd3149001301950464;
assign f1_rom[442] = 52'd3144603255439360;
assign f1_rom[443] = 52'd3144603255439360;
assign f1_rom[444] = 52'd3140205208928256;
assign f1_rom[445] = 52'd3140205208928256;
assign f1_rom[446] = 52'd3135807162417152;
assign f1_rom[447] = 52'd3135807162417152;
assign f1_rom[448] = 52'd3131409115906048;
assign f1_rom[449] = 52'd3131409115906048;
assign f1_rom[450] = 52'd3127011069394944;
assign f1_rom[451] = 52'd3127011069394944;
assign f1_rom[452] = 52'd3122613022883840;
assign f1_rom[453] = 52'd3122613022883840;
assign f1_rom[454] = 52'd3118214976372736;
assign f1_rom[455] = 52'd3118214976372736;
assign f1_rom[456] = 52'd3113816929861632;
assign f1_rom[457] = 52'd3113816929861632;
assign f1_rom[458] = 52'd3113816929861632;
assign f1_rom[459] = 52'd3109418883350528;
assign f1_rom[460] = 52'd3109418883350528;
assign f1_rom[461] = 52'd3105020836839424;
assign f1_rom[462] = 52'd3105020836839424;
assign f1_rom[463] = 52'd3100622790328320;
assign f1_rom[464] = 52'd3100622790328320;
assign f1_rom[465] = 52'd3096224743817216;
assign f1_rom[466] = 52'd3096224743817216;
assign f1_rom[467] = 52'd3091826697306112;
assign f1_rom[468] = 52'd3091826697306112;
assign f1_rom[469] = 52'd3087428650795008;
assign f1_rom[470] = 52'd3087428650795008;
assign f1_rom[471] = 52'd3083030604283904;
assign f1_rom[472] = 52'd3083030604283904;
assign f1_rom[473] = 52'd3078632557772800;
assign f1_rom[474] = 52'd3078632557772800;
assign f1_rom[475] = 52'd3078632557772800;
assign f1_rom[476] = 52'd3074234511261696;
assign f1_rom[477] = 52'd3074234511261696;
assign f1_rom[478] = 52'd3069836464750592;
assign f1_rom[479] = 52'd3069836464750592;
assign f1_rom[480] = 52'd3065438418239488;
assign f1_rom[481] = 52'd3065438418239488;
assign f1_rom[482] = 52'd3061040371728384;
assign f1_rom[483] = 52'd3061040371728384;
assign f1_rom[484] = 52'd3056642325217280;
assign f1_rom[485] = 52'd3056642325217280;
assign f1_rom[486] = 52'd3052244278706176;
assign f1_rom[487] = 52'd3052244278706176;
assign f1_rom[488] = 52'd3052244278706176;
assign f1_rom[489] = 52'd3047846232195072;
assign f1_rom[490] = 52'd3047846232195072;
assign f1_rom[491] = 52'd3043448185683968;
assign f1_rom[492] = 52'd3043448185683968;
assign f1_rom[493] = 52'd3039050139172864;
assign f1_rom[494] = 52'd3039050139172864;
assign f1_rom[495] = 52'd3034652092661760;
assign f1_rom[496] = 52'd3034652092661760;
assign f1_rom[497] = 52'd3030254046150656;
assign f1_rom[498] = 52'd3030254046150656;
assign f1_rom[499] = 52'd3025855999639552;
assign f1_rom[500] = 52'd3025855999639552;
assign f1_rom[501] = 52'd3025855999639552;
assign f1_rom[502] = 52'd3021457953128448;
assign f1_rom[503] = 52'd3021457953128448;
assign f1_rom[504] = 52'd3017059906617344;
assign f1_rom[505] = 52'd3017059906617344;
assign f1_rom[506] = 52'd3012661860106240;
assign f1_rom[507] = 52'd3012661860106240;
assign f1_rom[508] = 52'd3008263813595136;
assign f1_rom[509] = 52'd3008263813595136;
assign f1_rom[510] = 52'd3008263813595136;
assign f1_rom[511] = 52'd3003865767084032;
assign f1_rom[512] = 52'd3003865767084032;
assign f1_rom[513] = 52'd2999467720572928;
assign f1_rom[514] = 52'd2999467720572928;
assign f1_rom[515] = 52'd2995069674061824;
assign f1_rom[516] = 52'd2995069674061824;
assign f1_rom[517] = 52'd2990671627550720;
assign f1_rom[518] = 52'd2990671627550720;
assign f1_rom[519] = 52'd2990671627550720;
assign f1_rom[520] = 52'd2986273581039616;
assign f1_rom[521] = 52'd2986273581039616;
assign f1_rom[522] = 52'd2981875534528512;
assign f1_rom[523] = 52'd2981875534528512;
assign f1_rom[524] = 52'd2977477488017408;
assign f1_rom[525] = 52'd2977477488017408;
assign f1_rom[526] = 52'd2977477488017408;
assign f1_rom[527] = 52'd2973079441506304;
assign f1_rom[528] = 52'd2973079441506304;
assign f1_rom[529] = 52'd2968681394995200;
assign f1_rom[530] = 52'd2968681394995200;
assign f1_rom[531] = 52'd2964283348484096;
assign f1_rom[532] = 52'd2964283348484096;
assign f1_rom[533] = 52'd2959885301972992;
assign f1_rom[534] = 52'd2959885301972992;
assign f1_rom[535] = 52'd2959885301972992;
assign f1_rom[536] = 52'd2955487255461888;
assign f1_rom[537] = 52'd2955487255461888;
assign f1_rom[538] = 52'd2951089208950784;
assign f1_rom[539] = 52'd2951089208950784;
assign f1_rom[540] = 52'd2946691162439680;
assign f1_rom[541] = 52'd2946691162439680;
assign f1_rom[542] = 52'd2946691162439680;
assign f1_rom[543] = 52'd2942293115928576;
assign f1_rom[544] = 52'd2942293115928576;
assign f1_rom[545] = 52'd2937895069417472;
assign f1_rom[546] = 52'd2937895069417472;
assign f1_rom[547] = 52'd2933497022906368;
assign f1_rom[548] = 52'd2933497022906368;
assign f1_rom[549] = 52'd2933497022906368;
assign f1_rom[550] = 52'd2929098976395264;
assign f1_rom[551] = 52'd2929098976395264;
assign f1_rom[552] = 52'd2924700929884160;
assign f1_rom[553] = 52'd2924700929884160;
assign f1_rom[554] = 52'd2920302883373056;
assign f1_rom[555] = 52'd2920302883373056;
assign f1_rom[556] = 52'd2920302883373056;
assign f1_rom[557] = 52'd2915904836861952;
assign f1_rom[558] = 52'd2915904836861952;
assign f1_rom[559] = 52'd2911506790350848;
assign f1_rom[560] = 52'd2911506790350848;
assign f1_rom[561] = 52'd2911506790350848;
assign f1_rom[562] = 52'd2907108743839744;
assign f1_rom[563] = 52'd2907108743839744;
assign f1_rom[564] = 52'd2902710697328640;
assign f1_rom[565] = 52'd2902710697328640;
assign f1_rom[566] = 52'd2898312650817536;
assign f1_rom[567] = 52'd2898312650817536;
assign f1_rom[568] = 52'd2898312650817536;
assign f1_rom[569] = 52'd2893914604306432;
assign f1_rom[570] = 52'd2893914604306432;
assign f1_rom[571] = 52'd2889516557795328;
assign f1_rom[572] = 52'd2889516557795328;
assign f1_rom[573] = 52'd2889516557795328;
assign f1_rom[574] = 52'd2885118511284224;
assign f1_rom[575] = 52'd2885118511284224;
assign f1_rom[576] = 52'd2880720464773120;
assign f1_rom[577] = 52'd2880720464773120;
assign f1_rom[578] = 52'd2880720464773120;
assign f1_rom[579] = 52'd2876322418262016;
assign f1_rom[580] = 52'd2876322418262016;
assign f1_rom[581] = 52'd2871924371750912;
assign f1_rom[582] = 52'd2871924371750912;
assign f1_rom[583] = 52'd2871924371750912;
assign f1_rom[584] = 52'd2867526325239808;
assign f1_rom[585] = 52'd2867526325239808;
assign f1_rom[586] = 52'd2863128278728704;
assign f1_rom[587] = 52'd2863128278728704;
assign f1_rom[588] = 52'd2858730232217600;
assign f1_rom[589] = 52'd2858730232217600;
assign f1_rom[590] = 52'd2858730232217600;
assign f1_rom[591] = 52'd2854332185706496;
assign f1_rom[592] = 52'd2854332185706496;
assign f1_rom[593] = 52'd2849934139195392;
assign f1_rom[594] = 52'd2849934139195392;
assign f1_rom[595] = 52'd2849934139195392;
assign f1_rom[596] = 52'd2845536092684288;
assign f1_rom[597] = 52'd2845536092684288;
assign f1_rom[598] = 52'd2841138046173184;
assign f1_rom[599] = 52'd2841138046173184;
assign f1_rom[600] = 52'd2841138046173184;
assign f1_rom[601] = 52'd2836739999662080;
assign f1_rom[602] = 52'd2836739999662080;
assign f1_rom[603] = 52'd2832341953150976;
assign f1_rom[604] = 52'd2832341953150976;
assign f1_rom[605] = 52'd2832341953150976;
assign f1_rom[606] = 52'd2827943906639872;
assign f1_rom[607] = 52'd2827943906639872;
assign f1_rom[608] = 52'd2827943906639872;
assign f1_rom[609] = 52'd2823545860128768;
assign f1_rom[610] = 52'd2823545860128768;
assign f1_rom[611] = 52'd2819147813617664;
assign f1_rom[612] = 52'd2819147813617664;
assign f1_rom[613] = 52'd2819147813617664;
assign f1_rom[614] = 52'd2814749767106560;
assign f1_rom[615] = 52'd2814749767106560;
assign f1_rom[616] = 52'd2810351720595456;
assign f1_rom[617] = 52'd2810351720595456;
assign f1_rom[618] = 52'd2810351720595456;
assign f1_rom[619] = 52'd2805953674084352;
assign f1_rom[620] = 52'd2805953674084352;
assign f1_rom[621] = 52'd2801555627573248;
assign f1_rom[622] = 52'd2801555627573248;
assign f1_rom[623] = 52'd2801555627573248;
assign f1_rom[624] = 52'd2797157581062144;
assign f1_rom[625] = 52'd2797157581062144;
assign f1_rom[626] = 52'd2797157581062144;
assign f1_rom[627] = 52'd2792759534551040;
assign f1_rom[628] = 52'd2792759534551040;
assign f1_rom[629] = 52'd2788361488039936;
assign f1_rom[630] = 52'd2788361488039936;
assign f1_rom[631] = 52'd2788361488039936;
assign f1_rom[632] = 52'd2783963441528832;
assign f1_rom[633] = 52'd2783963441528832;
assign f1_rom[634] = 52'd2779565395017728;
assign f1_rom[635] = 52'd2779565395017728;
assign f1_rom[636] = 52'd2779565395017728;
assign f1_rom[637] = 52'd2775167348506624;
assign f1_rom[638] = 52'd2775167348506624;
assign f1_rom[639] = 52'd2775167348506624;
assign f1_rom[640] = 52'd2770769301995520;
assign f1_rom[641] = 52'd2770769301995520;
assign f1_rom[642] = 52'd2766371255484416;
assign f1_rom[643] = 52'd2766371255484416;
assign f1_rom[644] = 52'd2766371255484416;
assign f1_rom[645] = 52'd2761973208973312;
assign f1_rom[646] = 52'd2761973208973312;
assign f1_rom[647] = 52'd2761973208973312;
assign f1_rom[648] = 52'd2757575162462208;
assign f1_rom[649] = 52'd2757575162462208;
assign f1_rom[650] = 52'd2753177115951104;
assign f1_rom[651] = 52'd2753177115951104;
assign f1_rom[652] = 52'd2753177115951104;
assign f1_rom[653] = 52'd2748779069440000;
assign f1_rom[654] = 52'd2748779069440000;
assign f1_rom[655] = 52'd2748779069440000;
assign f1_rom[656] = 52'd2744381022928896;
assign f1_rom[657] = 52'd2744381022928896;
assign f1_rom[658] = 52'd2739982976417792;
assign f1_rom[659] = 52'd2739982976417792;
assign f1_rom[660] = 52'd2739982976417792;
assign f1_rom[661] = 52'd2735584929906688;
assign f1_rom[662] = 52'd2735584929906688;
assign f1_rom[663] = 52'd2735584929906688;
assign f1_rom[664] = 52'd2731186883395584;
assign f1_rom[665] = 52'd2731186883395584;
assign f1_rom[666] = 52'd2726788836884480;
assign f1_rom[667] = 52'd2726788836884480;
assign f1_rom[668] = 52'd2726788836884480;
assign f1_rom[669] = 52'd2722390790373376;
assign f1_rom[670] = 52'd2722390790373376;
assign f1_rom[671] = 52'd2722390790373376;
assign f1_rom[672] = 52'd2717992743862272;
assign f1_rom[673] = 52'd2717992743862272;
assign f1_rom[674] = 52'd2717992743862272;
assign f1_rom[675] = 52'd2713594697351168;
assign f1_rom[676] = 52'd2713594697351168;
assign f1_rom[677] = 52'd2709196650840064;
assign f1_rom[678] = 52'd2709196650840064;
assign f1_rom[679] = 52'd2709196650840064;
assign f1_rom[680] = 52'd2704798604328960;
assign f1_rom[681] = 52'd2704798604328960;
assign f1_rom[682] = 52'd2704798604328960;
assign f1_rom[683] = 52'd2700400557817856;
assign f1_rom[684] = 52'd2700400557817856;
assign f1_rom[685] = 52'd2700400557817856;
assign f1_rom[686] = 52'd2696002511306752;
assign f1_rom[687] = 52'd2696002511306752;
assign f1_rom[688] = 52'd2691604464795648;
assign f1_rom[689] = 52'd2691604464795648;
assign f1_rom[690] = 52'd2691604464795648;
assign f1_rom[691] = 52'd2687206418284544;
assign f1_rom[692] = 52'd2687206418284544;
assign f1_rom[693] = 52'd2687206418284544;
assign f1_rom[694] = 52'd2682808371773440;
assign f1_rom[695] = 52'd2682808371773440;
assign f1_rom[696] = 52'd2682808371773440;
assign f1_rom[697] = 52'd2678410325262336;
assign f1_rom[698] = 52'd2678410325262336;
assign f1_rom[699] = 52'd2678410325262336;
assign f1_rom[700] = 52'd2674012278751232;
assign f1_rom[701] = 52'd2674012278751232;
assign f1_rom[702] = 52'd2674012278751232;
assign f1_rom[703] = 52'd2669614232240128;
assign f1_rom[704] = 52'd2669614232240128;
assign f1_rom[705] = 52'd2665216185729024;
assign f1_rom[706] = 52'd2665216185729024;
assign f1_rom[707] = 52'd2665216185729024;
assign f1_rom[708] = 52'd2660818139217920;
assign f1_rom[709] = 52'd2660818139217920;
assign f1_rom[710] = 52'd2660818139217920;
assign f1_rom[711] = 52'd2656420092706816;
assign f1_rom[712] = 52'd2656420092706816;
assign f1_rom[713] = 52'd2656420092706816;
assign f1_rom[714] = 52'd2652022046195712;
assign f1_rom[715] = 52'd2652022046195712;
assign f1_rom[716] = 52'd2652022046195712;
assign f1_rom[717] = 52'd2647623999684608;
assign f1_rom[718] = 52'd2647623999684608;
assign f1_rom[719] = 52'd2647623999684608;
assign f1_rom[720] = 52'd2643225953173504;
assign f1_rom[721] = 52'd2643225953173504;
assign f1_rom[722] = 52'd2643225953173504;
assign f1_rom[723] = 52'd2638827906662400;
assign f1_rom[724] = 52'd2638827906662400;
assign f1_rom[725] = 52'd2638827906662400;
assign f1_rom[726] = 52'd2634429860151296;
assign f1_rom[727] = 52'd2634429860151296;
assign f1_rom[728] = 52'd2634429860151296;
assign f1_rom[729] = 52'd2630031813640192;
assign f1_rom[730] = 52'd2630031813640192;
assign f1_rom[731] = 52'd2625633767129088;
assign f1_rom[732] = 52'd2625633767129088;
assign f1_rom[733] = 52'd2625633767129088;
assign f1_rom[734] = 52'd2621235720617984;
assign f1_rom[735] = 52'd2621235720617984;
assign f1_rom[736] = 52'd2621235720617984;
assign f1_rom[737] = 52'd2616837674106880;
assign f1_rom[738] = 52'd2616837674106880;
assign f1_rom[739] = 52'd2616837674106880;
assign f1_rom[740] = 52'd2612439627595776;
assign f1_rom[741] = 52'd2612439627595776;
assign f1_rom[742] = 52'd2612439627595776;
assign f1_rom[743] = 52'd2608041581084672;
assign f1_rom[744] = 52'd2608041581084672;
assign f1_rom[745] = 52'd2608041581084672;
assign f1_rom[746] = 52'd2603643534573568;
assign f1_rom[747] = 52'd2603643534573568;
assign f1_rom[748] = 52'd2603643534573568;
assign f1_rom[749] = 52'd2599245488062464;
assign f1_rom[750] = 52'd2599245488062464;
assign f1_rom[751] = 52'd2599245488062464;
assign f1_rom[752] = 52'd2594847441551360;
assign f1_rom[753] = 52'd2594847441551360;
assign f1_rom[754] = 52'd2594847441551360;
assign f1_rom[755] = 52'd2590449395040256;
assign f1_rom[756] = 52'd2590449395040256;
assign f1_rom[757] = 52'd2590449395040256;
assign f1_rom[758] = 52'd2586051348529152;
assign f1_rom[759] = 52'd2586051348529152;
assign f1_rom[760] = 52'd2586051348529152;
assign f1_rom[761] = 52'd2581653302018048;
assign f1_rom[762] = 52'd2581653302018048;
assign f1_rom[763] = 52'd2581653302018048;
assign f1_rom[764] = 52'd2577255255506944;
assign f1_rom[765] = 52'd2577255255506944;
assign f1_rom[766] = 52'd2577255255506944;
assign f1_rom[767] = 52'd2572857208995840;
assign f1_rom[768] = 52'd2572857208995840;
assign f1_rom[769] = 52'd2572857208995840;
assign f1_rom[770] = 52'd2568459162484736;
assign f1_rom[771] = 52'd2568459162484736;
assign f1_rom[772] = 52'd2568459162484736;
assign f1_rom[773] = 52'd2568459162484736;
assign f1_rom[774] = 52'd2564061115973632;
assign f1_rom[775] = 52'd2564061115973632;
assign f1_rom[776] = 52'd2564061115973632;
assign f1_rom[777] = 52'd2559663069462528;
assign f1_rom[778] = 52'd2559663069462528;
assign f1_rom[779] = 52'd2559663069462528;
assign f1_rom[780] = 52'd2555265022951424;
assign f1_rom[781] = 52'd2555265022951424;
assign f1_rom[782] = 52'd2555265022951424;
assign f1_rom[783] = 52'd2550866976440320;
assign f1_rom[784] = 52'd2550866976440320;
assign f1_rom[785] = 52'd2550866976440320;
assign f1_rom[786] = 52'd2546468929929216;
assign f1_rom[787] = 52'd2546468929929216;
assign f1_rom[788] = 52'd2546468929929216;
assign f1_rom[789] = 52'd2542070883418112;
assign f1_rom[790] = 52'd2542070883418112;
assign f1_rom[791] = 52'd2542070883418112;
assign f1_rom[792] = 52'd2537672836907008;
assign f1_rom[793] = 52'd2537672836907008;
assign f1_rom[794] = 52'd2537672836907008;
assign f1_rom[795] = 52'd2533274790395904;
assign f1_rom[796] = 52'd2533274790395904;
assign f1_rom[797] = 52'd2533274790395904;
assign f1_rom[798] = 52'd2533274790395904;
assign f1_rom[799] = 52'd2528876743884800;
assign f1_rom[800] = 52'd2528876743884800;
assign f1_rom[801] = 52'd2528876743884800;
assign f1_rom[802] = 52'd2524478697373696;
assign f1_rom[803] = 52'd2524478697373696;
assign f1_rom[804] = 52'd2524478697373696;
assign f1_rom[805] = 52'd2520080650862592;
assign f1_rom[806] = 52'd2520080650862592;
assign f1_rom[807] = 52'd2520080650862592;
assign f1_rom[808] = 52'd2515682604351488;
assign f1_rom[809] = 52'd2515682604351488;
assign f1_rom[810] = 52'd2515682604351488;
assign f1_rom[811] = 52'd2511284557840384;
assign f1_rom[812] = 52'd2511284557840384;
assign f1_rom[813] = 52'd2511284557840384;
assign f1_rom[814] = 52'd2506886511329280;
assign f1_rom[815] = 52'd2506886511329280;
assign f1_rom[816] = 52'd2506886511329280;
assign f1_rom[817] = 52'd2506886511329280;
assign f1_rom[818] = 52'd2502488464818176;
assign f1_rom[819] = 52'd2502488464818176;
assign f1_rom[820] = 52'd2502488464818176;
assign f1_rom[821] = 52'd2498090418307072;
assign f1_rom[822] = 52'd2498090418307072;
assign f1_rom[823] = 52'd2498090418307072;
assign f1_rom[824] = 52'd2493692371795968;
assign f1_rom[825] = 52'd2493692371795968;
assign f1_rom[826] = 52'd2493692371795968;
assign f1_rom[827] = 52'd2489294325284864;
assign f1_rom[828] = 52'd2489294325284864;
assign f1_rom[829] = 52'd2489294325284864;
assign f1_rom[830] = 52'd2489294325284864;
assign f1_rom[831] = 52'd2484896278773760;
assign f1_rom[832] = 52'd2484896278773760;
assign f1_rom[833] = 52'd2484896278773760;
assign f1_rom[834] = 52'd2480498232262656;
assign f1_rom[835] = 52'd2480498232262656;
assign f1_rom[836] = 52'd2480498232262656;
assign f1_rom[837] = 52'd2476100185751552;
assign f1_rom[838] = 52'd2476100185751552;
assign f1_rom[839] = 52'd2476100185751552;
assign f1_rom[840] = 52'd2476100185751552;
assign f1_rom[841] = 52'd2471702139240448;
assign f1_rom[842] = 52'd2471702139240448;
assign f1_rom[843] = 52'd2471702139240448;
assign f1_rom[844] = 52'd2467304092729344;
assign f1_rom[845] = 52'd2467304092729344;
assign f1_rom[846] = 52'd2467304092729344;
assign f1_rom[847] = 52'd2462906046218240;
assign f1_rom[848] = 52'd2462906046218240;
assign f1_rom[849] = 52'd2462906046218240;
assign f1_rom[850] = 52'd2462906046218240;
assign f1_rom[851] = 52'd2458507999707136;
assign f1_rom[852] = 52'd2458507999707136;
assign f1_rom[853] = 52'd2458507999707136;
assign f1_rom[854] = 52'd2454109953196032;
assign f1_rom[855] = 52'd2454109953196032;
assign f1_rom[856] = 52'd2454109953196032;
assign f1_rom[857] = 52'd2449711906684928;
assign f1_rom[858] = 52'd2449711906684928;
assign f1_rom[859] = 52'd2449711906684928;
assign f1_rom[860] = 52'd2449711906684928;
assign f1_rom[861] = 52'd2445313860173824;
assign f1_rom[862] = 52'd2445313860173824;
assign f1_rom[863] = 52'd2445313860173824;
assign f1_rom[864] = 52'd2440915813662720;
assign f1_rom[865] = 52'd2440915813662720;
assign f1_rom[866] = 52'd2440915813662720;
assign f1_rom[867] = 52'd2440915813662720;
assign f1_rom[868] = 52'd2436517767151616;
assign f1_rom[869] = 52'd2436517767151616;
assign f1_rom[870] = 52'd2436517767151616;
assign f1_rom[871] = 52'd2432119720640512;
assign f1_rom[872] = 52'd2432119720640512;
assign f1_rom[873] = 52'd2432119720640512;
assign f1_rom[874] = 52'd2427721674129408;
assign f1_rom[875] = 52'd2427721674129408;
assign f1_rom[876] = 52'd2427721674129408;
assign f1_rom[877] = 52'd2427721674129408;
assign f1_rom[878] = 52'd2423323627618304;
assign f1_rom[879] = 52'd2423323627618304;
assign f1_rom[880] = 52'd2423323627618304;
assign f1_rom[881] = 52'd2418925581107200;
assign f1_rom[882] = 52'd2418925581107200;
assign f1_rom[883] = 52'd2418925581107200;
assign f1_rom[884] = 52'd2418925581107200;
assign f1_rom[885] = 52'd2414527534596096;
assign f1_rom[886] = 52'd2414527534596096;
assign f1_rom[887] = 52'd2414527534596096;
assign f1_rom[888] = 52'd2410129488084992;
assign f1_rom[889] = 52'd2410129488084992;
assign f1_rom[890] = 52'd2410129488084992;
assign f1_rom[891] = 52'd2410129488084992;
assign f1_rom[892] = 52'd2405731441573888;
assign f1_rom[893] = 52'd2405731441573888;
assign f1_rom[894] = 52'd2405731441573888;
assign f1_rom[895] = 52'd2401333395062784;
assign f1_rom[896] = 52'd2401333395062784;
assign f1_rom[897] = 52'd2401333395062784;
assign f1_rom[898] = 52'd2401333395062784;
assign f1_rom[899] = 52'd2396935348551680;
assign f1_rom[900] = 52'd2396935348551680;
assign f1_rom[901] = 52'd2396935348551680;
assign f1_rom[902] = 52'd2392537302040576;
assign f1_rom[903] = 52'd2392537302040576;
assign f1_rom[904] = 52'd2392537302040576;
assign f1_rom[905] = 52'd2392537302040576;
assign f1_rom[906] = 52'd2388139255529472;
assign f1_rom[907] = 52'd2388139255529472;
assign f1_rom[908] = 52'd2388139255529472;
assign f1_rom[909] = 52'd2383741209018368;
assign f1_rom[910] = 52'd2383741209018368;
assign f1_rom[911] = 52'd2383741209018368;
assign f1_rom[912] = 52'd2383741209018368;
assign f1_rom[913] = 52'd2379343162507264;
assign f1_rom[914] = 52'd2379343162507264;
assign f1_rom[915] = 52'd2379343162507264;
assign f1_rom[916] = 52'd2379343162507264;
assign f1_rom[917] = 52'd2374945115996160;
assign f1_rom[918] = 52'd2374945115996160;
assign f1_rom[919] = 52'd2374945115996160;
assign f1_rom[920] = 52'd2370547069485056;
assign f1_rom[921] = 52'd2370547069485056;
assign f1_rom[922] = 52'd2370547069485056;
assign f1_rom[923] = 52'd2370547069485056;
assign f1_rom[924] = 52'd2366149022973952;
assign f1_rom[925] = 52'd2366149022973952;
assign f1_rom[926] = 52'd2366149022973952;
assign f1_rom[927] = 52'd2361750976462848;
assign f1_rom[928] = 52'd2361750976462848;
assign f1_rom[929] = 52'd2361750976462848;
assign f1_rom[930] = 52'd2361750976462848;
assign f1_rom[931] = 52'd2357352929951744;
assign f1_rom[932] = 52'd2357352929951744;
assign f1_rom[933] = 52'd2357352929951744;
assign f1_rom[934] = 52'd2357352929951744;
assign f1_rom[935] = 52'd2352954883440640;
assign f1_rom[936] = 52'd2352954883440640;
assign f1_rom[937] = 52'd2352954883440640;
assign f1_rom[938] = 52'd2348556836929536;
assign f1_rom[939] = 52'd2348556836929536;
assign f1_rom[940] = 52'd2348556836929536;
assign f1_rom[941] = 52'd2348556836929536;
assign f1_rom[942] = 52'd2344158790418432;
assign f1_rom[943] = 52'd2344158790418432;
assign f1_rom[944] = 52'd2344158790418432;
assign f1_rom[945] = 52'd2344158790418432;
assign f1_rom[946] = 52'd2339760743907328;
assign f1_rom[947] = 52'd2339760743907328;
assign f1_rom[948] = 52'd2339760743907328;
assign f1_rom[949] = 52'd2335362697396224;
assign f1_rom[950] = 52'd2335362697396224;
assign f1_rom[951] = 52'd2335362697396224;
assign f1_rom[952] = 52'd2335362697396224;
assign f1_rom[953] = 52'd2330964650885120;
assign f1_rom[954] = 52'd2330964650885120;
assign f1_rom[955] = 52'd2330964650885120;
assign f1_rom[956] = 52'd2330964650885120;
assign f1_rom[957] = 52'd2326566604374016;
assign f1_rom[958] = 52'd2326566604374016;
assign f1_rom[959] = 52'd2326566604374016;
assign f1_rom[960] = 52'd2326566604374016;
assign f1_rom[961] = 52'd2322168557862912;
assign f1_rom[962] = 52'd2322168557862912;
assign f1_rom[963] = 52'd2322168557862912;
assign f1_rom[964] = 52'd2317770511351808;
assign f1_rom[965] = 52'd2317770511351808;
assign f1_rom[966] = 52'd2317770511351808;
assign f1_rom[967] = 52'd2317770511351808;
assign f1_rom[968] = 52'd2313372464840704;
assign f1_rom[969] = 52'd2313372464840704;
assign f1_rom[970] = 52'd2313372464840704;
assign f1_rom[971] = 52'd2313372464840704;
assign f1_rom[972] = 52'd2308974418329600;
assign f1_rom[973] = 52'd2308974418329600;
assign f1_rom[974] = 52'd2308974418329600;
assign f1_rom[975] = 52'd2308974418329600;
assign f1_rom[976] = 52'd2304576371818496;
assign f1_rom[977] = 52'd2304576371818496;
assign f1_rom[978] = 52'd2304576371818496;
assign f1_rom[979] = 52'd2304576371818496;
assign f1_rom[980] = 52'd2300178325307392;
assign f1_rom[981] = 52'd2300178325307392;
assign f1_rom[982] = 52'd2300178325307392;
assign f1_rom[983] = 52'd2295780278796288;
assign f1_rom[984] = 52'd2295780278796288;
assign f1_rom[985] = 52'd2295780278796288;
assign f1_rom[986] = 52'd2295780278796288;
assign f1_rom[987] = 52'd2291382232285184;
assign f1_rom[988] = 52'd2291382232285184;
assign f1_rom[989] = 52'd2291382232285184;
assign f1_rom[990] = 52'd2291382232285184;
assign f1_rom[991] = 52'd2286984185774080;
assign f1_rom[992] = 52'd2286984185774080;
assign f1_rom[993] = 52'd2286984185774080;
assign f1_rom[994] = 52'd2286984185774080;
assign f1_rom[995] = 52'd2282586139262976;
assign f1_rom[996] = 52'd2282586139262976;
assign f1_rom[997] = 52'd2282586139262976;
assign f1_rom[998] = 52'd2282586139262976;
assign f1_rom[999] = 52'd2278188092751872;
assign f1_rom[1000] = 52'd2278188092751872;
assign f1_rom[1001] = 52'd2278188092751872;
assign f1_rom[1002] = 52'd2278188092751872;
assign f1_rom[1003] = 52'd2273790046240768;
assign f1_rom[1004] = 52'd2273790046240768;
assign f1_rom[1005] = 52'd2273790046240768;
assign f1_rom[1006] = 52'd2273790046240768;
assign f1_rom[1007] = 52'd2269391999729664;
assign f1_rom[1008] = 52'd2269391999729664;
assign f1_rom[1009] = 52'd2269391999729664;
assign f1_rom[1010] = 52'd2269391999729664;
assign f1_rom[1011] = 52'd2264993953218560;
assign f1_rom[1012] = 52'd2264993953218560;
assign f1_rom[1013] = 52'd2264993953218560;
assign f1_rom[1014] = 52'd2264993953218560;
assign f1_rom[1015] = 52'd2260595906707456;
assign f1_rom[1016] = 52'd2260595906707456;
assign f1_rom[1017] = 52'd2260595906707456;
assign f1_rom[1018] = 52'd2260595906707456;
assign f1_rom[1019] = 52'd2256197860196352;
assign f1_rom[1020] = 52'd2256197860196352;
assign f1_rom[1021] = 52'd2256197860196352;
assign f1_rom[1022] = 52'd2256197860196352;
assign f1_rom[1023] = 52'd2251799813685248;

wire [51:0] f1_ln_rom [1023:0];
assign f1_ln_rom[0] = 52'd0;
assign f1_ln_rom[1] = 52'd4400195393878;  
assign f1_ln_rom[2] = 52'd8804694158020;  
assign f1_ln_rom[3] = 52'd13213504718019; 
assign f1_ln_rom[4] = 52'd17626635524235; 
assign f1_ln_rom[5] = 52'd22044095051897; 
assign f1_ln_rom[6] = 52'd26465891801195; 
assign f1_ln_rom[7] = 52'd30892034297384; 
assign f1_ln_rom[8] = 52'd35322531090877; 
assign f1_ln_rom[9] = 52'd39757390757348; 
assign f1_ln_rom[10] = 52'd44196621897830;
assign f1_ln_rom[11] = 52'd48640233138816;
assign f1_ln_rom[12] = 52'd53088233132357;
assign f1_ln_rom[13] = 52'd57540630556169;
assign f1_ln_rom[14] = 52'd61997434113726;
assign f1_ln_rom[15] = 52'd66458652534370;
assign f1_ln_rom[16] = 52'd70924294573409;
assign f1_ln_rom[17] = 52'd75394369012222;
assign f1_ln_rom[18] = 52'd79868884658361;
assign f1_ln_rom[19] = 52'd84347850345657;
assign f1_ln_rom[20] = 52'd88831274934323;
assign f1_ln_rom[21] = 52'd93319167311062;
assign f1_ln_rom[22] = 52'd97811536389167;
assign f1_ln_rom[23] = 52'd97811536389167;
assign f1_ln_rom[24] = 52'd102308391108635;
assign f1_ln_rom[25] = 52'd106809740436267;
assign f1_ln_rom[26] = 52'd111315593365778;
assign f1_ln_rom[27] = 52'd115825958917905;
assign f1_ln_rom[28] = 52'd120340846140516;
assign f1_ln_rom[29] = 52'd124860264108716;
assign f1_ln_rom[30] = 52'd129384221924960;
assign f1_ln_rom[31] = 52'd133912728719161;
assign f1_ln_rom[32] = 52'd138445793648801;
assign f1_ln_rom[33] = 52'd142983425899042;
assign f1_ln_rom[34] = 52'd147525634682837;
assign f1_ln_rom[35] = 52'd152072429241044;
assign f1_ln_rom[36] = 52'd156623818842538;
assign f1_ln_rom[37] = 52'd161179812784322;
assign f1_ln_rom[38] = 52'd165740420391645;
assign f1_ln_rom[39] = 52'd170305651018115;
assign f1_ln_rom[40] = 52'd170305651018115;
assign f1_ln_rom[41] = 52'd174875514045813;
assign f1_ln_rom[42] = 52'd179450018885407;
assign f1_ln_rom[43] = 52'd184029174976275;
assign f1_ln_rom[44] = 52'd188612991786615;
assign f1_ln_rom[45] = 52'd193201478813566;
assign f1_ln_rom[46] = 52'd197794645583323;
assign f1_ln_rom[47] = 52'd202392501651260;
assign f1_ln_rom[48] = 52'd206995056602046;
assign f1_ln_rom[49] = 52'd211602320049766;
assign f1_ln_rom[50] = 52'd216214301638042;
assign f1_ln_rom[51] = 52'd220831011040153;
assign f1_ln_rom[52] = 52'd220831011040153;
assign f1_ln_rom[53] = 52'd225452457959156;
assign f1_ln_rom[54] = 52'd230078652128012;
assign f1_ln_rom[55] = 52'd234709603309704;
assign f1_ln_rom[56] = 52'd239345321297365;
assign f1_ln_rom[57] = 52'd243985815914401;
assign f1_ln_rom[58] = 52'd248631097014613;
assign f1_ln_rom[59] = 52'd253281174482326;
assign f1_ln_rom[60] = 52'd257936058232515;
assign f1_ln_rom[61] = 52'd262595758210930;
assign f1_ln_rom[62] = 52'd262595758210930;
assign f1_ln_rom[63] = 52'd267260284394225;
assign f1_ln_rom[64] = 52'd271929646790084;
assign f1_ln_rom[65] = 52'd276603855437353;
assign f1_ln_rom[66] = 52'd281282920406168;
assign f1_ln_rom[67] = 52'd285966851798084;
assign f1_ln_rom[68] = 52'd290655659746208;
assign f1_ln_rom[69] = 52'd295349354415329;
assign f1_ln_rom[70] = 52'd300047946002051;
assign f1_ln_rom[71] = 52'd300047946002051;
assign f1_ln_rom[72] = 52'd304751444734925;
assign f1_ln_rom[73] = 52'd309459860874582;
assign f1_ln_rom[74] = 52'd314173204713873;
assign f1_ln_rom[75] = 52'd318891486577994;
assign f1_ln_rom[76] = 52'd323614716824631;
assign f1_ln_rom[77] = 52'd328342905844090;
assign f1_ln_rom[78] = 52'd328342905844090;
assign f1_ln_rom[79] = 52'd333076064059440;
assign f1_ln_rom[80] = 52'd337814201926645;
assign f1_ln_rom[81] = 52'd342557329934705;
assign f1_ln_rom[82] = 52'd347305458605798;
assign f1_ln_rom[83] = 52'd352058598495416;
assign f1_ln_rom[84] = 52'd356816760192507;
assign f1_ln_rom[85] = 52'd356816760192507;
assign f1_ln_rom[86] = 52'd361579954319618;
assign f1_ln_rom[87] = 52'd366348191533035;
assign f1_ln_rom[88] = 52'd371121482522929;
assign f1_ln_rom[89] = 52'd375899838013496;
assign f1_ln_rom[90] = 52'd380683268763106;
assign f1_ln_rom[91] = 52'd385471785564445;
assign f1_ln_rom[92] = 52'd385471785564445;
assign f1_ln_rom[93] = 52'd390265399244660;
assign f1_ln_rom[94] = 52'd395064120665512;
assign f1_ln_rom[95] = 52'd399867960723515;
assign f1_ln_rom[96] = 52'd404676930350094;
assign f1_ln_rom[97] = 52'd409491040511726;
assign f1_ln_rom[98] = 52'd409491040511726;
assign f1_ln_rom[99] = 52'd414310302210093;
assign f1_ln_rom[100] = 52'd419134726482237;
assign f1_ln_rom[101] = 52'd423964324400703;
assign f1_ln_rom[102] = 52'd428799107073700;
assign f1_ln_rom[103] = 52'd433639085645251;
assign f1_ln_rom[104] = 52'd433639085645251;
assign f1_ln_rom[105] = 52'd438484271295342;
assign f1_ln_rom[106] = 52'd443334675240089;
assign f1_ln_rom[107] = 52'd448190308731879;
assign f1_ln_rom[108] = 52'd453051183059540;
assign f1_ln_rom[109] = 52'd457917309548491;
assign f1_ln_rom[110] = 52'd457917309548491;
assign f1_ln_rom[111] = 52'd462788699560900;
assign f1_ln_rom[112] = 52'd467665364495846;
assign f1_ln_rom[113] = 52'd472547315789481;
assign f1_ln_rom[114] = 52'd477434564915184;
assign f1_ln_rom[115] = 52'd477434564915184;
assign f1_ln_rom[116] = 52'd482327123383730;
assign f1_ln_rom[117] = 52'd487225002743447;
assign f1_ln_rom[118] = 52'd492128214580385;
assign f1_ln_rom[119] = 52'd497036770518475;
assign f1_ln_rom[120] = 52'd497036770518475;
assign f1_ln_rom[121] = 52'd501950682219698;
assign f1_ln_rom[122] = 52'd506869961384250;
assign f1_ln_rom[123] = 52'd511794619750710;
assign f1_ln_rom[124] = 52'd516724669096206;
assign f1_ln_rom[125] = 52'd516724669096206;
assign f1_ln_rom[126] = 52'd521660121236586;
assign f1_ln_rom[127] = 52'd526600988026588;
assign f1_ln_rom[128] = 52'd531547281360008;
assign f1_ln_rom[129] = 52'd536499013169876;
assign f1_ln_rom[130] = 52'd536499013169876;
assign f1_ln_rom[131] = 52'd541456195428626;
assign f1_ln_rom[132] = 52'd546418840148270;
assign f1_ln_rom[133] = 52'd551386959380574;
assign f1_ln_rom[134] = 52'd551386959380574;
assign f1_ln_rom[135] = 52'd556360565217230;
assign f1_ln_rom[136] = 52'd561339669790038;
assign f1_ln_rom[137] = 52'd566324285271080;
assign f1_ln_rom[138] = 52'd571314423872898;
assign f1_ln_rom[139] = 52'd571314423872898;
assign f1_ln_rom[140] = 52'd576310097848675;
assign f1_ln_rom[141] = 52'd581311319492417;
assign f1_ln_rom[142] = 52'd586318101139131;
assign f1_ln_rom[143] = 52'd586318101139131;
assign f1_ln_rom[144] = 52'd591330455165010;
assign f1_ln_rom[145] = 52'd596348393987615;
assign f1_ln_rom[146] = 52'd601371930066064;
assign f1_ln_rom[147] = 52'd606401075901208;
assign f1_ln_rom[148] = 52'd606401075901208;
assign f1_ln_rom[149] = 52'd611435844035830;
assign f1_ln_rom[150] = 52'd616476247054822;
assign f1_ln_rom[151] = 52'd621522297585381;
assign f1_ln_rom[152] = 52'd621522297585381;
assign f1_ln_rom[153] = 52'd626574008297194;
assign f1_ln_rom[154] = 52'd631631391902632;
assign f1_ln_rom[155] = 52'd636694461156940;
assign f1_ln_rom[156] = 52'd636694461156940;
assign f1_ln_rom[157] = 52'd641763228858432;
assign f1_ln_rom[158] = 52'd646837707848683;
assign f1_ln_rom[159] = 52'd651917911012725;
assign f1_ln_rom[160] = 52'd651917911012725;
assign f1_ln_rom[161] = 52'd657003851279243;
assign f1_ln_rom[162] = 52'd662095541620775;
assign f1_ln_rom[163] = 52'd667192995053907;
assign f1_ln_rom[164] = 52'd667192995053907;
assign f1_ln_rom[165] = 52'd672296224639473;
assign f1_ln_rom[166] = 52'd677405243482758;
assign f1_ln_rom[167] = 52'd682520064733699;
assign f1_ln_rom[168] = 52'd682520064733699;
assign f1_ln_rom[169] = 52'd687640701587087;
assign f1_ln_rom[170] = 52'd692767167282773;
assign f1_ln_rom[171] = 52'd697899475105872;
assign f1_ln_rom[172] = 52'd697899475105872;
assign f1_ln_rom[173] = 52'd703037638386970;
assign f1_ln_rom[174] = 52'd708181670502330;
assign f1_ln_rom[175] = 52'd708181670502330;
assign f1_ln_rom[176] = 52'd713331584874108;
assign f1_ln_rom[177] = 52'd718487394970551;
assign f1_ln_rom[178] = 52'd723649114306220;
assign f1_ln_rom[179] = 52'd723649114306220;
assign f1_ln_rom[180] = 52'd728816756442196;
assign f1_ln_rom[181] = 52'd733990334986297;
assign f1_ln_rom[182] = 52'd739169863593289;
assign f1_ln_rom[183] = 52'd739169863593289;
assign f1_ln_rom[184] = 52'd744355355965106;
assign f1_ln_rom[185] = 52'd749546825851066;
assign f1_ln_rom[186] = 52'd749546825851066;
assign f1_ln_rom[187] = 52'd754744287048092;
assign f1_ln_rom[188] = 52'd759947753400926;
assign f1_ln_rom[189] = 52'd765157238802358;
assign f1_ln_rom[190] = 52'd765157238802358;
assign f1_ln_rom[191] = 52'd770372757193443;
assign f1_ln_rom[192] = 52'd775594322563727;
assign f1_ln_rom[193] = 52'd775594322563727;
assign f1_ln_rom[194] = 52'd780821948951471;
assign f1_ln_rom[195] = 52'd786055650443879;
assign f1_ln_rom[196] = 52'd791295441177326;
assign f1_ln_rom[197] = 52'd791295441177326;
assign f1_ln_rom[198] = 52'd796541335337584;
assign f1_ln_rom[199] = 52'd801793347160057;
assign f1_ln_rom[200] = 52'd801793347160057;
assign f1_ln_rom[201] = 52'd807051490930008;
assign f1_ln_rom[202] = 52'd812315780982794;
assign f1_ln_rom[203] = 52'd812315780982794;
assign f1_ln_rom[204] = 52'd817586231704106;
assign f1_ln_rom[205] = 52'd822862857530193;
assign f1_ln_rom[206] = 52'd822862857530193;
assign f1_ln_rom[207] = 52'd828145672948110;
assign f1_ln_rom[208] = 52'd833434692495954;
assign f1_ln_rom[209] = 52'd838729930763098;
assign f1_ln_rom[210] = 52'd838729930763098;
assign f1_ln_rom[211] = 52'd844031402390442;
assign f1_ln_rom[212] = 52'd849339122070648;
assign f1_ln_rom[213] = 52'd849339122070648;
assign f1_ln_rom[214] = 52'd854653104548390;
assign f1_ln_rom[215] = 52'd859973364620594;
assign f1_ln_rom[216] = 52'd859973364620594;
assign f1_ln_rom[217] = 52'd865299917136693;
assign f1_ln_rom[218] = 52'd870632776998866;
assign f1_ln_rom[219] = 52'd870632776998866;
assign f1_ln_rom[220] = 52'd875971959162296;
assign f1_ln_rom[221] = 52'd881317478635419;
assign f1_ln_rom[222] = 52'd881317478635419;
assign f1_ln_rom[223] = 52'd886669350480177;
assign f1_ln_rom[224] = 52'd892027589812272;
assign f1_ln_rom[225] = 52'd892027589812272;
assign f1_ln_rom[226] = 52'd897392211801423;
assign f1_ln_rom[227] = 52'd902763231671623;
assign f1_ln_rom[228] = 52'd902763231671623;
assign f1_ln_rom[229] = 52'd908140664701400;
assign f1_ln_rom[230] = 52'd913524526224076;
assign f1_ln_rom[231] = 52'd913524526224076;
assign f1_ln_rom[232] = 52'd918914831628030;
assign f1_ln_rom[233] = 52'd924311596356961;
assign f1_ln_rom[234] = 52'd924311596356961;
assign f1_ln_rom[235] = 52'd929714835910154;
assign f1_ln_rom[236] = 52'd935124565842748;
assign f1_ln_rom[237] = 52'd935124565842748;
assign f1_ln_rom[238] = 52'd940540801766006;
assign f1_ln_rom[239] = 52'd945963559347578;
assign f1_ln_rom[240] = 52'd945963559347578;
assign f1_ln_rom[241] = 52'd951392854311785;
assign f1_ln_rom[242] = 52'd956828702439880;
assign f1_ln_rom[243] = 52'd956828702439880;
assign f1_ln_rom[244] = 52'd962271119570331;
assign f1_ln_rom[245] = 52'd967720121599098;
assign f1_ln_rom[246] = 52'd967720121599098;
assign f1_ln_rom[247] = 52'd973175724479907;
assign f1_ln_rom[248] = 52'd978637944224534;
assign f1_ln_rom[249] = 52'd978637944224534;
assign f1_ln_rom[250] = 52'd984106796903084;
assign f1_ln_rom[251] = 52'd989582298644278;
assign f1_ln_rom[252] = 52'd989582298644278;
assign f1_ln_rom[253] = 52'd995064465635738;
assign f1_ln_rom[254] = 52'd1000553314124270;
assign f1_ln_rom[255] = 52'd1000553314124270;
assign f1_ln_rom[256] = 52'd1006048860416158;
assign f1_ln_rom[257] = 52'd1006048860416158;
assign f1_ln_rom[258] = 52'd1011551120877450;
assign f1_ln_rom[259] = 52'd1017060111934257;
assign f1_ln_rom[260] = 52'd1017060111934257;
assign f1_ln_rom[261] = 52'd1022575850073039;
assign f1_ln_rom[262] = 52'd1028098351840909;
assign f1_ln_rom[263] = 52'd1028098351840909;
assign f1_ln_rom[264] = 52'd1033627633845923;
assign f1_ln_rom[265] = 52'd1039163712757386;
assign f1_ln_rom[266] = 52'd1039163712757386;
assign f1_ln_rom[267] = 52'd1044706605306152;
assign f1_ln_rom[268] = 52'd1044706605306152;
assign f1_ln_rom[269] = 52'd1050256328284925;
assign f1_ln_rom[270] = 52'd1055812898548567;
assign f1_ln_rom[271] = 52'd1055812898548567;
assign f1_ln_rom[272] = 52'd1061376333014402;
assign f1_ln_rom[273] = 52'd1066946648662530;
assign f1_ln_rom[274] = 52'd1066946648662530;
assign f1_ln_rom[275] = 52'd1072523862536133;
assign f1_ln_rom[276] = 52'd1072523862536133;
assign f1_ln_rom[277] = 52'd1078107991741791;
assign f1_ln_rom[278] = 52'd1083699053449793;
assign f1_ln_rom[279] = 52'd1083699053449793;
assign f1_ln_rom[280] = 52'd1089297064894461;
assign f1_ln_rom[281] = 52'd1089297064894461;
assign f1_ln_rom[282] = 52'd1094902043374460;
assign f1_ln_rom[283] = 52'd1100514006253125;
assign f1_ln_rom[284] = 52'd1100514006253125;
assign f1_ln_rom[285] = 52'd1106132970958782;
assign f1_ln_rom[286] = 52'd1111758954985071;
assign f1_ln_rom[287] = 52'd1111758954985071;
assign f1_ln_rom[288] = 52'd1117391975891276;
assign f1_ln_rom[289] = 52'd1117391975891276;
assign f1_ln_rom[290] = 52'd1123032051302650;
assign f1_ln_rom[291] = 52'd1128679198910749;
assign f1_ln_rom[292] = 52'd1128679198910749;
assign f1_ln_rom[293] = 52'd1134333436473764;
assign f1_ln_rom[294] = 52'd1134333436473764;
assign f1_ln_rom[295] = 52'd1139994781816856;
assign f1_ln_rom[296] = 52'd1145663252832494;
assign f1_ln_rom[297] = 52'd1145663252832494;
assign f1_ln_rom[298] = 52'd1151338867480790;
assign f1_ln_rom[299] = 52'd1151338867480790;
assign f1_ln_rom[300] = 52'd1157021643789848;
assign f1_ln_rom[301] = 52'd1162711599856102;
assign f1_ln_rom[302] = 52'd1162711599856102;
assign f1_ln_rom[303] = 52'd1168408753844661;
assign f1_ln_rom[304] = 52'd1168408753844661;
assign f1_ln_rom[305] = 52'd1174113123989662;
assign f1_ln_rom[306] = 52'd1179824728594617;
assign f1_ln_rom[307] = 52'd1179824728594617;
assign f1_ln_rom[308] = 52'd1185543586032764;
assign f1_ln_rom[309] = 52'd1185543586032764;
assign f1_ln_rom[310] = 52'd1191269714747424;
assign f1_ln_rom[311] = 52'd1197003133252359;
assign f1_ln_rom[312] = 52'd1197003133252359;
assign f1_ln_rom[313] = 52'd1202743860132127;
assign f1_ln_rom[314] = 52'd1202743860132127;
assign f1_ln_rom[315] = 52'd1208491914042447;
assign f1_ln_rom[316] = 52'd1208491914042447;
assign f1_ln_rom[317] = 52'd1214247313710561;
assign f1_ln_rom[318] = 52'd1220010077935601;
assign f1_ln_rom[319] = 52'd1220010077935601;
assign f1_ln_rom[320] = 52'd1225780225588957;
assign f1_ln_rom[321] = 52'd1225780225588957;
assign f1_ln_rom[322] = 52'd1231557775614648;
assign f1_ln_rom[323] = 52'd1237342747029694;
assign f1_ln_rom[324] = 52'd1237342747029694;
assign f1_ln_rom[325] = 52'd1243135158924496;
assign f1_ln_rom[326] = 52'd1243135158924496;
assign f1_ln_rom[327] = 52'd1248935030463205;
assign f1_ln_rom[328] = 52'd1248935030463205;
assign f1_ln_rom[329] = 52'd1254742380884113;
assign f1_ln_rom[330] = 52'd1260557229500029;
assign f1_ln_rom[331] = 52'd1260557229500029;
assign f1_ln_rom[332] = 52'd1266379595698666;
assign f1_ln_rom[333] = 52'd1266379595698666;
assign f1_ln_rom[334] = 52'd1272209498943029;
assign f1_ln_rom[335] = 52'd1272209498943029;
assign f1_ln_rom[336] = 52'd1278046958771807;
assign f1_ln_rom[337] = 52'd1283891994799762;
assign f1_ln_rom[338] = 52'd1283891994799762;
assign f1_ln_rom[339] = 52'd1289744626718130;
assign f1_ln_rom[340] = 52'd1289744626718130;
assign f1_ln_rom[341] = 52'd1295604874295012;
assign f1_ln_rom[342] = 52'd1295604874295012;
assign f1_ln_rom[343] = 52'd1301472757375783;
assign f1_ln_rom[344] = 52'd1301472757375783;
assign f1_ln_rom[345] = 52'd1307348295883487;
assign f1_ln_rom[346] = 52'd1313231509819248;
assign f1_ln_rom[347] = 52'd1313231509819248;
assign f1_ln_rom[348] = 52'd1319122419262677;
assign f1_ln_rom[349] = 52'd1319122419262677;
assign f1_ln_rom[350] = 52'd1325021044372284;
assign f1_ln_rom[351] = 52'd1325021044372284;
assign f1_ln_rom[352] = 52'd1330927405385890;
assign f1_ln_rom[353] = 52'd1336841522621045;
assign f1_ln_rom[354] = 52'd1336841522621045;
assign f1_ln_rom[355] = 52'd1342763416475449;
assign f1_ln_rom[356] = 52'd1342763416475449;
assign f1_ln_rom[357] = 52'd1348693107427370;
assign f1_ln_rom[358] = 52'd1348693107427370;
assign f1_ln_rom[359] = 52'd1354630616036072;
assign f1_ln_rom[360] = 52'd1354630616036072;
assign f1_ln_rom[361] = 52'd1360575962942243;
assign f1_ln_rom[362] = 52'd1360575962942243;
assign f1_ln_rom[363] = 52'd1366529168868422;
assign f1_ln_rom[364] = 52'd1372490254619436;
assign f1_ln_rom[365] = 52'd1372490254619436;
assign f1_ln_rom[366] = 52'd1378459241082837;
assign f1_ln_rom[367] = 52'd1378459241082837;
assign f1_ln_rom[368] = 52'd1384436149229336;
assign f1_ln_rom[369] = 52'd1384436149229336;
assign f1_ln_rom[370] = 52'd1390421000113249;
assign f1_ln_rom[371] = 52'd1390421000113249;
assign f1_ln_rom[372] = 52'd1396413814872942;
assign f1_ln_rom[373] = 52'd1396413814872942;
assign f1_ln_rom[374] = 52'd1402414614731280;
assign f1_ln_rom[375] = 52'd1402414614731280;
assign f1_ln_rom[376] = 52'd1408423420996071;
assign f1_ln_rom[377] = 52'd1414440255060530;
assign f1_ln_rom[378] = 52'd1414440255060530;
assign f1_ln_rom[379] = 52'd1420465138403728;
assign f1_ln_rom[380] = 52'd1420465138403728;
assign f1_ln_rom[381] = 52'd1426498092591058;
assign f1_ln_rom[382] = 52'd1426498092591058;
assign f1_ln_rom[383] = 52'd1432539139274693;
assign f1_ln_rom[384] = 52'd1432539139274693;
assign f1_ln_rom[385] = 52'd1438588300194055;
assign f1_ln_rom[386] = 52'd1438588300194055;
assign f1_ln_rom[387] = 52'd1444645597176284;
assign f1_ln_rom[388] = 52'd1444645597176284;
assign f1_ln_rom[389] = 52'd1450711052136712;
assign f1_ln_rom[390] = 52'd1450711052136712;
assign f1_ln_rom[391] = 52'd1456784687079334;
assign f1_ln_rom[392] = 52'd1456784687079334;
assign f1_ln_rom[393] = 52'd1462866524097295;
assign f1_ln_rom[394] = 52'd1468956585373362;
assign f1_ln_rom[395] = 52'd1468956585373362;
assign f1_ln_rom[396] = 52'd1475054893180420;
assign f1_ln_rom[397] = 52'd1475054893180420;
assign f1_ln_rom[398] = 52'd1481161469881951;
assign f1_ln_rom[399] = 52'd1481161469881951;
assign f1_ln_rom[400] = 52'd1487276337932534;
assign f1_ln_rom[401] = 52'd1487276337932534;
assign f1_ln_rom[402] = 52'd1493399519878336;
assign f1_ln_rom[403] = 52'd1493399519878336;
assign f1_ln_rom[404] = 52'd1499531038357610;
assign f1_ln_rom[405] = 52'd1499531038357610;
assign f1_ln_rom[406] = 52'd1505670916101203;
assign f1_ln_rom[407] = 52'd1505670916101203;
assign f1_ln_rom[408] = 52'd1511819175933055;
assign f1_ln_rom[409] = 52'd1511819175933055;
assign f1_ln_rom[410] = 52'd1517975840770710;
assign f1_ln_rom[411] = 52'd1517975840770710;
assign f1_ln_rom[412] = 52'd1524140933625832;
assign f1_ln_rom[413] = 52'd1524140933625832;
assign f1_ln_rom[414] = 52'd1530314477604716;
assign f1_ln_rom[415] = 52'd1530314477604716;
assign f1_ln_rom[416] = 52'd1536496495908812;
assign f1_ln_rom[417] = 52'd1536496495908812;
assign f1_ln_rom[418] = 52'd1542687011835244;
assign f1_ln_rom[419] = 52'd1542687011835244;
assign f1_ln_rom[420] = 52'd1548886048777339;
assign f1_ln_rom[421] = 52'd1548886048777339;
assign f1_ln_rom[422] = 52'd1555093630225160;
assign f1_ln_rom[423] = 52'd1555093630225160;
assign f1_ln_rom[424] = 52'd1561309779766034;
assign f1_ln_rom[425] = 52'd1561309779766034;
assign f1_ln_rom[426] = 52'd1567534521085096;
assign f1_ln_rom[427] = 52'd1567534521085096;
assign f1_ln_rom[428] = 52'd1573767877965827;
assign f1_ln_rom[429] = 52'd1573767877965827;
assign f1_ln_rom[430] = 52'd1580009874290597;
assign f1_ln_rom[431] = 52'd1580009874290597;
assign f1_ln_rom[432] = 52'd1586260534041221;
assign f1_ln_rom[433] = 52'd1586260534041221;
assign f1_ln_rom[434] = 52'd1592519881299505;
assign f1_ln_rom[435] = 52'd1592519881299505;
assign f1_ln_rom[436] = 52'd1598787940247807;
assign f1_ln_rom[437] = 52'd1598787940247807;
assign f1_ln_rom[438] = 52'd1605064735169595;
assign f1_ln_rom[439] = 52'd1605064735169595;
assign f1_ln_rom[440] = 52'd1611350290450012;
assign f1_ln_rom[441] = 52'd1611350290450012;
assign f1_ln_rom[442] = 52'd1617644630576447;
assign f1_ln_rom[443] = 52'd1617644630576447;
assign f1_ln_rom[444] = 52'd1623947780139103;
assign f1_ln_rom[445] = 52'd1623947780139103;
assign f1_ln_rom[446] = 52'd1630259763831576;
assign f1_ln_rom[447] = 52'd1630259763831576;
assign f1_ln_rom[448] = 52'd1636580606451436;
assign f1_ln_rom[449] = 52'd1636580606451436;
assign f1_ln_rom[450] = 52'd1642910332900811;
assign f1_ln_rom[451] = 52'd1642910332900811;
assign f1_ln_rom[452] = 52'd1649248968186973;
assign f1_ln_rom[453] = 52'd1649248968186973;
assign f1_ln_rom[454] = 52'd1655596537422936;
assign f1_ln_rom[455] = 52'd1655596537422936;
assign f1_ln_rom[456] = 52'd1661953065828048;
assign f1_ln_rom[457] = 52'd1661953065828048;
assign f1_ln_rom[458] = 52'd1661953065828048;
assign f1_ln_rom[459] = 52'd1668318578728594;
assign f1_ln_rom[460] = 52'd1668318578728594;
assign f1_ln_rom[461] = 52'd1674693101558404;
assign f1_ln_rom[462] = 52'd1674693101558404;
assign f1_ln_rom[463] = 52'd1681076659859457;
assign f1_ln_rom[464] = 52'd1681076659859457;
assign f1_ln_rom[465] = 52'd1687469279282503;
assign f1_ln_rom[466] = 52'd1687469279282503;
assign f1_ln_rom[467] = 52'd1693870985587673;
assign f1_ln_rom[468] = 52'd1693870985587673;
assign f1_ln_rom[469] = 52'd1700281804645107;
assign f1_ln_rom[470] = 52'd1700281804645107;
assign f1_ln_rom[471] = 52'd1706701762435580;
assign f1_ln_rom[472] = 52'd1706701762435580;
assign f1_ln_rom[473] = 52'd1713130885051135;
assign f1_ln_rom[474] = 52'd1713130885051135;
assign f1_ln_rom[475] = 52'd1713130885051135;
assign f1_ln_rom[476] = 52'd1719569198695716;
assign f1_ln_rom[477] = 52'd1719569198695716;
assign f1_ln_rom[478] = 52'd1726016729685812;
assign f1_ln_rom[479] = 52'd1726016729685812;
assign f1_ln_rom[480] = 52'd1732473504451101;
assign f1_ln_rom[481] = 52'd1732473504451101;
assign f1_ln_rom[482] = 52'd1738939549535101;
assign f1_ln_rom[483] = 52'd1738939549535101;
assign f1_ln_rom[484] = 52'd1745414891595824;
assign f1_ln_rom[485] = 52'd1745414891595824;
assign f1_ln_rom[486] = 52'd1751899557406433;
assign f1_ln_rom[487] = 52'd1751899557406433;
assign f1_ln_rom[488] = 52'd1751899557406433;
assign f1_ln_rom[489] = 52'd1758393573855912;
assign f1_ln_rom[490] = 52'd1758393573855912;
assign f1_ln_rom[491] = 52'd1764896967949730;
assign f1_ln_rom[492] = 52'd1764896967949730;
assign f1_ln_rom[493] = 52'd1771409766810518;
assign f1_ln_rom[494] = 52'd1771409766810518;
assign f1_ln_rom[495] = 52'd1777931997678742;
assign f1_ln_rom[496] = 52'd1777931997678742;
assign f1_ln_rom[497] = 52'd1784463687913397;
assign f1_ln_rom[498] = 52'd1784463687913397;
assign f1_ln_rom[499] = 52'd1791004864992684;
assign f1_ln_rom[500] = 52'd1791004864992684;
assign f1_ln_rom[501] = 52'd1791004864992684;
assign f1_ln_rom[502] = 52'd1797555556514711;
assign f1_ln_rom[503] = 52'd1797555556514711;
assign f1_ln_rom[504] = 52'd1804115790198190;
assign f1_ln_rom[505] = 52'd1804115790198190;
assign f1_ln_rom[506] = 52'd1810685593883141;
assign f1_ln_rom[507] = 52'd1810685593883141;
assign f1_ln_rom[508] = 52'd1817264995531599;
assign f1_ln_rom[509] = 52'd1817264995531599;
assign f1_ln_rom[510] = 52'd1817264995531599;
assign f1_ln_rom[511] = 52'd1823854023228328;
assign f1_ln_rom[512] = 52'd1823854023228328;
assign f1_ln_rom[513] = 52'd1830452705181545;
assign f1_ln_rom[514] = 52'd1830452705181545;
assign f1_ln_rom[515] = 52'd1837061069723638;
assign f1_ln_rom[516] = 52'd1837061069723638;
assign f1_ln_rom[517] = 52'd1843679145311902;
assign f1_ln_rom[518] = 52'd1843679145311902;
assign f1_ln_rom[519] = 52'd1843679145311902;
assign f1_ln_rom[520] = 52'd1850306960529269;
assign f1_ln_rom[521] = 52'd1850306960529269;
assign f1_ln_rom[522] = 52'd1856944544085051;
assign f1_ln_rom[523] = 52'd1856944544085051;
assign f1_ln_rom[524] = 52'd1863591924815688;
assign f1_ln_rom[525] = 52'd1863591924815688;
assign f1_ln_rom[526] = 52'd1863591924815688;
assign f1_ln_rom[527] = 52'd1870249131685497;
assign f1_ln_rom[528] = 52'd1870249131685497;
assign f1_ln_rom[529] = 52'd1876916193787430;
assign f1_ln_rom[530] = 52'd1876916193787430;
assign f1_ln_rom[531] = 52'd1883593140343836;
assign f1_ln_rom[532] = 52'd1883593140343836;
assign f1_ln_rom[533] = 52'd1890280000707232;
assign f1_ln_rom[534] = 52'd1890280000707232;
assign f1_ln_rom[535] = 52'd1890280000707232;
assign f1_ln_rom[536] = 52'd1896976804361076;
assign f1_ln_rom[537] = 52'd1896976804361076;
assign f1_ln_rom[538] = 52'd1903683580920545;
assign f1_ln_rom[539] = 52'd1903683580920545;
assign f1_ln_rom[540] = 52'd1910400360133324;
assign f1_ln_rom[541] = 52'd1910400360133324;
assign f1_ln_rom[542] = 52'd1910400360133324;
assign f1_ln_rom[543] = 52'd1917127171880394;
assign f1_ln_rom[544] = 52'd1917127171880394;
assign f1_ln_rom[545] = 52'd1923864046176834;
assign f1_ln_rom[546] = 52'd1923864046176834;
assign f1_ln_rom[547] = 52'd1930611013172622;
assign f1_ln_rom[548] = 52'd1930611013172622;
assign f1_ln_rom[549] = 52'd1930611013172622;
assign f1_ln_rom[550] = 52'd1937368103153445;
assign f1_ln_rom[551] = 52'd1937368103153445;
assign f1_ln_rom[552] = 52'd1944135346541512;
assign f1_ln_rom[553] = 52'd1944135346541512;
assign f1_ln_rom[554] = 52'd1950912773896383;
assign f1_ln_rom[555] = 52'd1950912773896383;
assign f1_ln_rom[556] = 52'd1950912773896383;
assign f1_ln_rom[557] = 52'd1957700415915788;
assign f1_ln_rom[558] = 52'd1957700415915788;
assign f1_ln_rom[559] = 52'd1964498303436468;
assign f1_ln_rom[560] = 52'd1964498303436468;
assign f1_ln_rom[561] = 52'd1964498303436468;
assign f1_ln_rom[562] = 52'd1971306467435014;
assign f1_ln_rom[563] = 52'd1971306467435014;
assign f1_ln_rom[564] = 52'd1978124939028712;
assign f1_ln_rom[565] = 52'd1978124939028712;
assign f1_ln_rom[566] = 52'd1984953749476396;
assign f1_ln_rom[567] = 52'd1984953749476396;
assign f1_ln_rom[568] = 52'd1984953749476396;
assign f1_ln_rom[569] = 52'd1991792930179312;
assign f1_ln_rom[570] = 52'd1991792930179312;
assign f1_ln_rom[571] = 52'd1998642512681982;
assign f1_ln_rom[572] = 52'd1998642512681982;
assign f1_ln_rom[573] = 52'd1998642512681982;
assign f1_ln_rom[574] = 52'd2005502528673074;
assign f1_ln_rom[575] = 52'd2005502528673074;
assign f1_ln_rom[576] = 52'd2012373009986287;
assign f1_ln_rom[577] = 52'd2012373009986287;
assign f1_ln_rom[578] = 52'd2012373009986287;
assign f1_ln_rom[579] = 52'd2019253988601233;
assign f1_ln_rom[580] = 52'd2019253988601233;
assign f1_ln_rom[581] = 52'd2026145496644332;
assign f1_ln_rom[582] = 52'd2026145496644332;
assign f1_ln_rom[583] = 52'd2026145496644332;
assign f1_ln_rom[584] = 52'd2033047566389713;
assign f1_ln_rom[585] = 52'd2033047566389713;
assign f1_ln_rom[586] = 52'd2039960230260118;
assign f1_ln_rom[587] = 52'd2039960230260118;
assign f1_ln_rom[588] = 52'd2046883520827820;
assign f1_ln_rom[589] = 52'd2046883520827820;
assign f1_ln_rom[590] = 52'd2046883520827820;
assign f1_ln_rom[591] = 52'd2053817470815538;
assign f1_ln_rom[592] = 52'd2053817470815538;
assign f1_ln_rom[593] = 52'd2060762113097371;
assign f1_ln_rom[594] = 52'd2060762113097371;
assign f1_ln_rom[595] = 52'd2060762113097371;
assign f1_ln_rom[596] = 52'd2067717480699730;
assign f1_ln_rom[597] = 52'd2067717480699730;
assign f1_ln_rom[598] = 52'd2074683606802280;
assign f1_ln_rom[599] = 52'd2074683606802280;
assign f1_ln_rom[600] = 52'd2074683606802280;
assign f1_ln_rom[601] = 52'd2081660524738892;
assign f1_ln_rom[602] = 52'd2081660524738892;
assign f1_ln_rom[603] = 52'd2088648267998598;
assign f1_ln_rom[604] = 52'd2088648267998598;
assign f1_ln_rom[605] = 52'd2088648267998598;
assign f1_ln_rom[606] = 52'd2095646870226555;
assign f1_ln_rom[607] = 52'd2095646870226555;
assign f1_ln_rom[608] = 52'd2095646870226555;
assign f1_ln_rom[609] = 52'd2102656365225020;
assign f1_ln_rom[610] = 52'd2102656365225020;
assign f1_ln_rom[611] = 52'd2109676786954327;
assign f1_ln_rom[612] = 52'd2109676786954327;
assign f1_ln_rom[613] = 52'd2109676786954327;
assign f1_ln_rom[614] = 52'd2116708169533876;
assign f1_ln_rom[615] = 52'd2116708169533876;
assign f1_ln_rom[616] = 52'd2123750547243123;
assign f1_ln_rom[617] = 52'd2123750547243123;
assign f1_ln_rom[618] = 52'd2123750547243123;
assign f1_ln_rom[619] = 52'd2130803954522592;
assign f1_ln_rom[620] = 52'd2130803954522592;
assign f1_ln_rom[621] = 52'd2137868425974876;
assign f1_ln_rom[622] = 52'd2137868425974876;
assign f1_ln_rom[623] = 52'd2137868425974876;
assign f1_ln_rom[624] = 52'd2144943996365661;
assign f1_ln_rom[625] = 52'd2144943996365661;
assign f1_ln_rom[626] = 52'd2144943996365661;
assign f1_ln_rom[627] = 52'd2152030700624752;
assign f1_ln_rom[628] = 52'd2152030700624752;
assign f1_ln_rom[629] = 52'd2159128573847107;
assign f1_ln_rom[630] = 52'd2159128573847107;
assign f1_ln_rom[631] = 52'd2159128573847107;
assign f1_ln_rom[632] = 52'd2166237651293878;
assign f1_ln_rom[633] = 52'd2166237651293878;
assign f1_ln_rom[634] = 52'd2173357968393465;
assign f1_ln_rom[635] = 52'd2173357968393465;
assign f1_ln_rom[636] = 52'd2173357968393465;
assign f1_ln_rom[637] = 52'd2180489560742574;
assign f1_ln_rom[638] = 52'd2180489560742574;
assign f1_ln_rom[639] = 52'd2180489560742574;
assign f1_ln_rom[640] = 52'd2187632464107284;
assign f1_ln_rom[641] = 52'd2187632464107284;
assign f1_ln_rom[642] = 52'd2194786714424126;
assign f1_ln_rom[643] = 52'd2194786714424126;
assign f1_ln_rom[644] = 52'd2194786714424126;
assign f1_ln_rom[645] = 52'd2201952347801163;
assign f1_ln_rom[646] = 52'd2201952347801163;
assign f1_ln_rom[647] = 52'd2201952347801163;
assign f1_ln_rom[648] = 52'd2209129400519089;
assign f1_ln_rom[649] = 52'd2209129400519089;
assign f1_ln_rom[650] = 52'd2216317909032327;
assign f1_ln_rom[651] = 52'd2216317909032327;
assign f1_ln_rom[652] = 52'd2216317909032327;
assign f1_ln_rom[653] = 52'd2223517909970142;
assign f1_ln_rom[654] = 52'd2223517909970142;
assign f1_ln_rom[655] = 52'd2223517909970142;
assign f1_ln_rom[656] = 52'd2230729440137761;
assign f1_ln_rom[657] = 52'd2230729440137761;
assign f1_ln_rom[658] = 52'd2237952536517500;
assign f1_ln_rom[659] = 52'd2237952536517500;
assign f1_ln_rom[660] = 52'd2237952536517500;
assign f1_ln_rom[661] = 52'd2245187236269904;
assign f1_ln_rom[662] = 52'd2245187236269904;
assign f1_ln_rom[663] = 52'd2245187236269904;
assign f1_ln_rom[664] = 52'd2252433576734892;
assign f1_ln_rom[665] = 52'd2252433576734892;
assign f1_ln_rom[666] = 52'd2259691595432918;
assign f1_ln_rom[667] = 52'd2259691595432918;
assign f1_ln_rom[668] = 52'd2259691595432918;
assign f1_ln_rom[669] = 52'd2266961330066128;
assign f1_ln_rom[670] = 52'd2266961330066128;
assign f1_ln_rom[671] = 52'd2266961330066128;
assign f1_ln_rom[672] = 52'd2274242818519546;
assign f1_ln_rom[673] = 52'd2274242818519546;
assign f1_ln_rom[674] = 52'd2274242818519546;
assign f1_ln_rom[675] = 52'd2281536098862249;
assign f1_ln_rom[676] = 52'd2281536098862249;
assign f1_ln_rom[677] = 52'd2288841209348566;
assign f1_ln_rom[678] = 52'd2288841209348566;
assign f1_ln_rom[679] = 52'd2288841209348566;
assign f1_ln_rom[680] = 52'd2296158188419282;
assign f1_ln_rom[681] = 52'd2296158188419282;
assign f1_ln_rom[682] = 52'd2296158188419282;
assign f1_ln_rom[683] = 52'd2303487074702851;
assign f1_ln_rom[684] = 52'd2303487074702851;
assign f1_ln_rom[685] = 52'd2303487074702851;
assign f1_ln_rom[686] = 52'd2310827907016617;
assign f1_ln_rom[687] = 52'd2310827907016617;
assign f1_ln_rom[688] = 52'd2318180724368052;
assign f1_ln_rom[689] = 52'd2318180724368052;
assign f1_ln_rom[690] = 52'd2318180724368052;
assign f1_ln_rom[691] = 52'd2325545565955998;
assign f1_ln_rom[692] = 52'd2325545565955998;
assign f1_ln_rom[693] = 52'd2325545565955998;
assign f1_ln_rom[694] = 52'd2332922471171918;
assign f1_ln_rom[695] = 52'd2332922471171918;
assign f1_ln_rom[696] = 52'd2332922471171918;
assign f1_ln_rom[697] = 52'd2340311479601164;
assign f1_ln_rom[698] = 52'd2340311479601164;
assign f1_ln_rom[699] = 52'd2340311479601164;
assign f1_ln_rom[700] = 52'd2347712631024253;
assign f1_ln_rom[701] = 52'd2347712631024253;
assign f1_ln_rom[702] = 52'd2347712631024253;
assign f1_ln_rom[703] = 52'd2355125965418144;
assign f1_ln_rom[704] = 52'd2355125965418144;
assign f1_ln_rom[705] = 52'd2362551522957543;
assign f1_ln_rom[706] = 52'd2362551522957543;
assign f1_ln_rom[707] = 52'd2362551522957543;
assign f1_ln_rom[708] = 52'd2369989344016202;
assign f1_ln_rom[709] = 52'd2369989344016202;
assign f1_ln_rom[710] = 52'd2369989344016202;
assign f1_ln_rom[711] = 52'd2377439469168240;
assign f1_ln_rom[712] = 52'd2377439469168240;
assign f1_ln_rom[713] = 52'd2377439469168240;
assign f1_ln_rom[714] = 52'd2384901939189474;
assign f1_ln_rom[715] = 52'd2384901939189474;
assign f1_ln_rom[716] = 52'd2384901939189474;
assign f1_ln_rom[717] = 52'd2392376795058747;
assign f1_ln_rom[718] = 52'd2392376795058747;
assign f1_ln_rom[719] = 52'd2392376795058747;
assign f1_ln_rom[720] = 52'd2399864077959292;
assign f1_ln_rom[721] = 52'd2399864077959292;
assign f1_ln_rom[722] = 52'd2399864077959292;
assign f1_ln_rom[723] = 52'd2407363829280084;
assign f1_ln_rom[724] = 52'd2407363829280084;
assign f1_ln_rom[725] = 52'd2407363829280084;
assign f1_ln_rom[726] = 52'd2414876090617216;
assign f1_ln_rom[727] = 52'd2414876090617216;
assign f1_ln_rom[728] = 52'd2414876090617216;
assign f1_ln_rom[729] = 52'd2422400903775282;
assign f1_ln_rom[730] = 52'd2422400903775282;
assign f1_ln_rom[731] = 52'd2429938310768777;
assign f1_ln_rom[732] = 52'd2429938310768777;
assign f1_ln_rom[733] = 52'd2429938310768777;
assign f1_ln_rom[734] = 52'd2437488353823497;
assign f1_ln_rom[735] = 52'd2437488353823497;
assign f1_ln_rom[736] = 52'd2437488353823497;
assign f1_ln_rom[737] = 52'd2445051075377966;
assign f1_ln_rom[738] = 52'd2445051075377966;
assign f1_ln_rom[739] = 52'd2445051075377966;
assign f1_ln_rom[740] = 52'd2452626518084861;
assign f1_ln_rom[741] = 52'd2452626518084861;
assign f1_ln_rom[742] = 52'd2452626518084861;
assign f1_ln_rom[743] = 52'd2460214724812462;
assign f1_ln_rom[744] = 52'd2460214724812462;
assign f1_ln_rom[745] = 52'd2460214724812462;
assign f1_ln_rom[746] = 52'd2467815738646099;
assign f1_ln_rom[747] = 52'd2467815738646099;
assign f1_ln_rom[748] = 52'd2467815738646099;
assign f1_ln_rom[749] = 52'd2475429602889630;
assign f1_ln_rom[750] = 52'd2475429602889630;
assign f1_ln_rom[751] = 52'd2475429602889630;
assign f1_ln_rom[752] = 52'd2483056361066910;
assign f1_ln_rom[753] = 52'd2483056361066910;
assign f1_ln_rom[754] = 52'd2483056361066910;
assign f1_ln_rom[755] = 52'd2490696056923296;
assign f1_ln_rom[756] = 52'd2490696056923296;
assign f1_ln_rom[757] = 52'd2490696056923296;
assign f1_ln_rom[758] = 52'd2498348734427140;
assign f1_ln_rom[759] = 52'd2498348734427140;
assign f1_ln_rom[760] = 52'd2498348734427140;
assign f1_ln_rom[761] = 52'd2506014437771318;
assign f1_ln_rom[762] = 52'd2506014437771318;
assign f1_ln_rom[763] = 52'd2506014437771318;
assign f1_ln_rom[764] = 52'd2513693211374754;
assign f1_ln_rom[765] = 52'd2513693211374754;
assign f1_ln_rom[766] = 52'd2513693211374754;
assign f1_ln_rom[767] = 52'd2521385099883970;
assign f1_ln_rom[768] = 52'd2521385099883970;
assign f1_ln_rom[769] = 52'd2521385099883970;
assign f1_ln_rom[770] = 52'd2529090148174636;
assign f1_ln_rom[771] = 52'd2529090148174636;
assign f1_ln_rom[772] = 52'd2529090148174636;
assign f1_ln_rom[773] = 52'd2529090148174636;
assign f1_ln_rom[774] = 52'd2536808401353151;
assign f1_ln_rom[775] = 52'd2536808401353151;
assign f1_ln_rom[776] = 52'd2536808401353151;
assign f1_ln_rom[777] = 52'd2544539904758218;
assign f1_ln_rom[778] = 52'd2544539904758218;
assign f1_ln_rom[779] = 52'd2544539904758218;
assign f1_ln_rom[780] = 52'd2552284703962446;
assign f1_ln_rom[781] = 52'd2552284703962446;
assign f1_ln_rom[782] = 52'd2552284703962446;
assign f1_ln_rom[783] = 52'd2560042844773964;
assign f1_ln_rom[784] = 52'd2560042844773964;
assign f1_ln_rom[785] = 52'd2560042844773964;
assign f1_ln_rom[786] = 52'd2567814373238042;
assign f1_ln_rom[787] = 52'd2567814373238042;
assign f1_ln_rom[788] = 52'd2567814373238042;
assign f1_ln_rom[789] = 52'd2575599335638733;
assign f1_ln_rom[790] = 52'd2575599335638733;
assign f1_ln_rom[791] = 52'd2575599335638733;
assign f1_ln_rom[792] = 52'd2583397778500529;
assign f1_ln_rom[793] = 52'd2583397778500529;
assign f1_ln_rom[794] = 52'd2583397778500529;
assign f1_ln_rom[795] = 52'd2591209748590025;
assign f1_ln_rom[796] = 52'd2591209748590025;
assign f1_ln_rom[797] = 52'd2591209748590025;
assign f1_ln_rom[798] = 52'd2591209748590025;
assign f1_ln_rom[799] = 52'd2599035292917605;
assign f1_ln_rom[800] = 52'd2599035292917605;
assign f1_ln_rom[801] = 52'd2599035292917605;
assign f1_ln_rom[802] = 52'd2606874458739138;
assign f1_ln_rom[803] = 52'd2606874458739138;
assign f1_ln_rom[804] = 52'd2606874458739138;
assign f1_ln_rom[805] = 52'd2614727293557690;
assign f1_ln_rom[806] = 52'd2614727293557690;
assign f1_ln_rom[807] = 52'd2614727293557690;
assign f1_ln_rom[808] = 52'd2622593845125252;
assign f1_ln_rom[809] = 52'd2622593845125252;
assign f1_ln_rom[810] = 52'd2622593845125252;
assign f1_ln_rom[811] = 52'd2630474161444482;
assign f1_ln_rom[812] = 52'd2630474161444482;
assign f1_ln_rom[813] = 52'd2630474161444482;
assign f1_ln_rom[814] = 52'd2638368290770462;
assign f1_ln_rom[815] = 52'd2638368290770462;
assign f1_ln_rom[816] = 52'd2638368290770462;
assign f1_ln_rom[817] = 52'd2638368290770462;
assign f1_ln_rom[818] = 52'd2646276281612472;
assign f1_ln_rom[819] = 52'd2646276281612472;
assign f1_ln_rom[820] = 52'd2646276281612472;
assign f1_ln_rom[821] = 52'd2654198182735778;
assign f1_ln_rom[822] = 52'd2654198182735778;
assign f1_ln_rom[823] = 52'd2654198182735778;
assign f1_ln_rom[824] = 52'd2662134043163434;
assign f1_ln_rom[825] = 52'd2662134043163434;
assign f1_ln_rom[826] = 52'd2662134043163434;
assign f1_ln_rom[827] = 52'd2670083912178109;
assign f1_ln_rom[828] = 52'd2670083912178109;
assign f1_ln_rom[829] = 52'd2670083912178109;
assign f1_ln_rom[830] = 52'd2670083912178109;
assign f1_ln_rom[831] = 52'd2678047839323914;
assign f1_ln_rom[832] = 52'd2678047839323914;
assign f1_ln_rom[833] = 52'd2678047839323914;
assign f1_ln_rom[834] = 52'd2686025874408262;
assign f1_ln_rom[835] = 52'd2686025874408262;
assign f1_ln_rom[836] = 52'd2686025874408262;
assign f1_ln_rom[837] = 52'd2694018067503733;
assign f1_ln_rom[838] = 52'd2694018067503733;
assign f1_ln_rom[839] = 52'd2694018067503733;
assign f1_ln_rom[840] = 52'd2694018067503733;
assign f1_ln_rom[841] = 52'd2702024468949963;
assign f1_ln_rom[842] = 52'd2702024468949963;
assign f1_ln_rom[843] = 52'd2702024468949963;
assign f1_ln_rom[844] = 52'd2710045129355542;
assign f1_ln_rom[845] = 52'd2710045129355542;
assign f1_ln_rom[846] = 52'd2710045129355542;
assign f1_ln_rom[847] = 52'd2718080099599939;
assign f1_ln_rom[848] = 52'd2718080099599939;
assign f1_ln_rom[849] = 52'd2718080099599939;
assign f1_ln_rom[850] = 52'd2718080099599939;
assign f1_ln_rom[851] = 52'd2726129430835432;
assign f1_ln_rom[852] = 52'd2726129430835432;
assign f1_ln_rom[853] = 52'd2726129430835432;
assign f1_ln_rom[854] = 52'd2734193174489068;
assign f1_ln_rom[855] = 52'd2734193174489068;
assign f1_ln_rom[856] = 52'd2734193174489068;
assign f1_ln_rom[857] = 52'd2742271382264629;
assign f1_ln_rom[858] = 52'd2742271382264629;
assign f1_ln_rom[859] = 52'd2742271382264629;
assign f1_ln_rom[860] = 52'd2742271382264629;
assign f1_ln_rom[861] = 52'd2750364106144628;
assign f1_ln_rom[862] = 52'd2750364106144628;
assign f1_ln_rom[863] = 52'd2750364106144628;
assign f1_ln_rom[864] = 52'd2758471398392308;
assign f1_ln_rom[865] = 52'd2758471398392308;
assign f1_ln_rom[866] = 52'd2758471398392308;
assign f1_ln_rom[867] = 52'd2758471398392308;
assign f1_ln_rom[868] = 52'd2766593311553672;
assign f1_ln_rom[869] = 52'd2766593311553672;
assign f1_ln_rom[870] = 52'd2766593311553672;
assign f1_ln_rom[871] = 52'd2774729898459528;
assign f1_ln_rom[872] = 52'd2774729898459528;
assign f1_ln_rom[873] = 52'd2774729898459528;
assign f1_ln_rom[874] = 52'd2782881212227546;
assign f1_ln_rom[875] = 52'd2782881212227546;
assign f1_ln_rom[876] = 52'd2782881212227546;
assign f1_ln_rom[877] = 52'd2782881212227546;
assign f1_ln_rom[878] = 52'd2791047306264342;
assign f1_ln_rom[879] = 52'd2791047306264342;
assign f1_ln_rom[880] = 52'd2791047306264342;
assign f1_ln_rom[881] = 52'd2799228234267574;
assign f1_ln_rom[882] = 52'd2799228234267574;
assign f1_ln_rom[883] = 52'd2799228234267574;
assign f1_ln_rom[884] = 52'd2799228234267574;
assign f1_ln_rom[885] = 52'd2807424050228068;
assign f1_ln_rom[886] = 52'd2807424050228068;
assign f1_ln_rom[887] = 52'd2807424050228068;
assign f1_ln_rom[888] = 52'd2815634808431946;
assign f1_ln_rom[889] = 52'd2815634808431946;
assign f1_ln_rom[890] = 52'd2815634808431946;
assign f1_ln_rom[891] = 52'd2815634808431946;
assign f1_ln_rom[892] = 52'd2823860563462792;
assign f1_ln_rom[893] = 52'd2823860563462792;
assign f1_ln_rom[894] = 52'd2823860563462792;
assign f1_ln_rom[895] = 52'd2832101370203824;
assign f1_ln_rom[896] = 52'd2832101370203824;
assign f1_ln_rom[897] = 52'd2832101370203824;
assign f1_ln_rom[898] = 52'd2832101370203824;
assign f1_ln_rom[899] = 52'd2840357283840096;
assign f1_ln_rom[900] = 52'd2840357283840096;
assign f1_ln_rom[901] = 52'd2840357283840096;
assign f1_ln_rom[902] = 52'd2848628359860706;
assign f1_ln_rom[903] = 52'd2848628359860706;
assign f1_ln_rom[904] = 52'd2848628359860706;
assign f1_ln_rom[905] = 52'd2848628359860706;
assign f1_ln_rom[906] = 52'd2856914654061047;
assign f1_ln_rom[907] = 52'd2856914654061047;
assign f1_ln_rom[908] = 52'd2856914654061047;
assign f1_ln_rom[909] = 52'd2865216222545053;
assign f1_ln_rom[910] = 52'd2865216222545053;
assign f1_ln_rom[911] = 52'd2865216222545053;
assign f1_ln_rom[912] = 52'd2865216222545053;
assign f1_ln_rom[913] = 52'd2873533121727486;
assign f1_ln_rom[914] = 52'd2873533121727486;
assign f1_ln_rom[915] = 52'd2873533121727486;
assign f1_ln_rom[916] = 52'd2873533121727486;
assign f1_ln_rom[917] = 52'd2881865408336234;
assign f1_ln_rom[918] = 52'd2881865408336234;
assign f1_ln_rom[919] = 52'd2881865408336234;
assign f1_ln_rom[920] = 52'd2890213139414630;
assign f1_ln_rom[921] = 52'd2890213139414630;
assign f1_ln_rom[922] = 52'd2890213139414630;
assign f1_ln_rom[923] = 52'd2890213139414630;
assign f1_ln_rom[924] = 52'd2898576372323800;
assign f1_ln_rom[925] = 52'd2898576372323800;
assign f1_ln_rom[926] = 52'd2898576372323800;
assign f1_ln_rom[927] = 52'd2906955164745025;
assign f1_ln_rom[928] = 52'd2906955164745025;
assign f1_ln_rom[929] = 52'd2906955164745025;
assign f1_ln_rom[930] = 52'd2906955164745025;
assign f1_ln_rom[931] = 52'd2915349574682128;
assign f1_ln_rom[932] = 52'd2915349574682128;
assign f1_ln_rom[933] = 52'd2915349574682128;
assign f1_ln_rom[934] = 52'd2915349574682128;
assign f1_ln_rom[935] = 52'd2923759660463883;
assign f1_ln_rom[936] = 52'd2923759660463883;
assign f1_ln_rom[937] = 52'd2923759660463883;
assign f1_ln_rom[938] = 52'd2932185480746449;
assign f1_ln_rom[939] = 52'd2932185480746449;
assign f1_ln_rom[940] = 52'd2932185480746449;
assign f1_ln_rom[941] = 52'd2932185480746449;
assign f1_ln_rom[942] = 52'd2940627094515822;
assign f1_ln_rom[943] = 52'd2940627094515822;
assign f1_ln_rom[944] = 52'd2940627094515822;
assign f1_ln_rom[945] = 52'd2940627094515822;
assign f1_ln_rom[946] = 52'd2949084561090316;
assign f1_ln_rom[947] = 52'd2949084561090316;
assign f1_ln_rom[948] = 52'd2949084561090316;
assign f1_ln_rom[949] = 52'd2957557940123060;
assign f1_ln_rom[950] = 52'd2957557940123060;
assign f1_ln_rom[951] = 52'd2957557940123060;
assign f1_ln_rom[952] = 52'd2957557940123060;
assign f1_ln_rom[953] = 52'd2966047291604524;
assign f1_ln_rom[954] = 52'd2966047291604524;
assign f1_ln_rom[955] = 52'd2966047291604524;
assign f1_ln_rom[956] = 52'd2966047291604524;
assign f1_ln_rom[957] = 52'd2974552675865068;
assign f1_ln_rom[958] = 52'd2974552675865068;
assign f1_ln_rom[959] = 52'd2974552675865068;
assign f1_ln_rom[960] = 52'd2974552675865068;
assign f1_ln_rom[961] = 52'd2983074153577516;
assign f1_ln_rom[962] = 52'd2983074153577516;
assign f1_ln_rom[963] = 52'd2983074153577516;
assign f1_ln_rom[964] = 52'd2991611785759748;
assign f1_ln_rom[965] = 52'd2991611785759748;
assign f1_ln_rom[966] = 52'd2991611785759748;
assign f1_ln_rom[967] = 52'd2991611785759748;
assign f1_ln_rom[968] = 52'd3000165633777329;
assign f1_ln_rom[969] = 52'd3000165633777329;
assign f1_ln_rom[970] = 52'd3000165633777329;
assign f1_ln_rom[971] = 52'd3000165633777329;
assign f1_ln_rom[972] = 52'd3008735759346148;
assign f1_ln_rom[973] = 52'd3008735759346148;
assign f1_ln_rom[974] = 52'd3008735759346148;
assign f1_ln_rom[975] = 52'd3008735759346148;
assign f1_ln_rom[976] = 52'd3017322224535091;
assign f1_ln_rom[977] = 52'd3017322224535091;
assign f1_ln_rom[978] = 52'd3017322224535091;
assign f1_ln_rom[979] = 52'd3017322224535091;
assign f1_ln_rom[980] = 52'd3025925091768746;
assign f1_ln_rom[981] = 52'd3025925091768746;
assign f1_ln_rom[982] = 52'd3025925091768746;
assign f1_ln_rom[983] = 52'd3034544423830114;
assign f1_ln_rom[984] = 52'd3034544423830114;
assign f1_ln_rom[985] = 52'd3034544423830114;
assign f1_ln_rom[986] = 52'd3034544423830114;
assign f1_ln_rom[987] = 52'd3043180283863368;
assign f1_ln_rom[988] = 52'd3043180283863368;
assign f1_ln_rom[989] = 52'd3043180283863368;
assign f1_ln_rom[990] = 52'd3043180283863368;
assign f1_ln_rom[991] = 52'd3051832735376624;
assign f1_ln_rom[992] = 52'd3051832735376624;
assign f1_ln_rom[993] = 52'd3051832735376624;
assign f1_ln_rom[994] = 52'd3051832735376624;
assign f1_ln_rom[995] = 52'd3060501842244743;
assign f1_ln_rom[996] = 52'd3060501842244743;
assign f1_ln_rom[997] = 52'd3060501842244743;
assign f1_ln_rom[998] = 52'd3060501842244743;
assign f1_ln_rom[999] = 52'd3069187668712162;
assign f1_ln_rom[1000] = 52'd3069187668712162;
assign f1_ln_rom[1001] = 52'd3069187668712162;
assign f1_ln_rom[1002] = 52'd3069187668712162;
assign f1_ln_rom[1003] = 52'd3077890279395752;
assign f1_ln_rom[1004] = 52'd3077890279395752;
assign f1_ln_rom[1005] = 52'd3077890279395752;
assign f1_ln_rom[1006] = 52'd3077890279395752;
assign f1_ln_rom[1007] = 52'd3086609739287696;
assign f1_ln_rom[1008] = 52'd3086609739287696;
assign f1_ln_rom[1009] = 52'd3086609739287696;
assign f1_ln_rom[1010] = 52'd3086609739287696;
assign f1_ln_rom[1011] = 52'd3095346113758409;
assign f1_ln_rom[1012] = 52'd3095346113758409;
assign f1_ln_rom[1013] = 52'd3095346113758409;
assign f1_ln_rom[1014] = 52'd3095346113758409;
assign f1_ln_rom[1015] = 52'd3104099468559474;
assign f1_ln_rom[1016] = 52'd3104099468559474;
assign f1_ln_rom[1017] = 52'd3104099468559474;
assign f1_ln_rom[1018] = 52'd3104099468559474;
assign f1_ln_rom[1019] = 52'd3112869869826612;
assign f1_ln_rom[1020] = 52'd3112869869826612;
assign f1_ln_rom[1021] = 52'd3112869869826612;
assign f1_ln_rom[1022] = 52'd3112869869826612;
assign f1_ln_rom[1023] = 52'd3121657384082680;

wire [10:0] shift;
wire shift_pn;

wire [52:0] f1;
wire [51:0] f1_ln;
wire [9:0] rom_index;

reg [10:0] shift_buffer [ITERATION_NUM-1:0];
reg shift_pn_buffer [ITERATION_NUM-1:0];
reg signed [52:0] f1_ln_buffer [ITERATION_NUM-1:0];

wire [52:0] x0;
wire [53+53-1:0] x1_full;
wire [52:0] x1;

//wire [22:0] ln;
wire signed [42:0] a;

//layer0
wire signed [42+42:0] layer0_value0_full; //a^2
reg signed [32:0] layer0_value0; 
reg signed [41:0] layer0_value1; // a/3
reg signed [42:0] a_buffer;

//layer1
reg signed [42:0] layer1_value0; //a-(a^2)/2
wire signed [32+32:0] layer1_value1_full; //a^2 * a^2
wire signed [41+32:0] layer1_value2_full; // (a^3)/3
reg signed [12:0] layer1_value1;
reg signed [21:0] layer1_value2;

//layer2 
reg signed [42:0] layer2_value0; //layer1_value0 - layer1_value1/4 + layer1_value2

wire in_NaN;
wire in_INF;
wire invalid_op;
wire overflow;
wire underflow;

reg invalid_op_buffer[ITERATION_NUM-1:0];
reg overflow_buffer[ITERATION_NUM-1:0];
reg in_valid_buffer[ITERATION_NUM-1:0];

wire [63:0] ln;
wire signed [53:0] ln_0;
wire [61:0] ln2_value;

wire    [5:0]   index;
wire    [31:0]   tmp4;
wire    [15:0]   tmp3;
wire    [7:0]   tmp0;
wire    [3:0]   tmp1;
wire    [1:0]   tmp2;
wire [63:0] ln_value;

wire [FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-1:0] ln_float0;

wire [63:0] ln_value_shift;

assign shift_pn = i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] >= 11'd1023 ? 0 : 1; 
assign shift = i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] >= 11'd1023 ? i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] - 1023 : 1023 - i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1];
 
assign rom_index = i_data[FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-11];
assign f1 = f1_rom[rom_index];
assign f1_ln = f1_ln_rom[rom_index];

assign x0 = {1'b1,i_data[FLOAT_FRAC_WIDTH-2:0]};
assign x1_full = (x0 * f1) >>> 52;
assign x1 = x1_full[52:0];

assign a = x1 - (1 <<< 52);

assign layer0_value0_full = a * a;

assign layer1_value1_full = layer0_value0 * layer0_value0;
assign layer1_value2_full = layer0_value0 * layer0_value1;

integer i0;
integer i1;
integer i2;
always @ ( posedge i_clk or negedge i_rst_n )
    if( !i_rst_n )
    begin
    for (i0 = 0; i0 < ITERATION_NUM; i0 = i0+1) begin
      shift_buffer[i0] <= 0;
      shift_pn_buffer[i0] <= 0;
      f1_ln_buffer[i0] <= 0;
    end
    
    layer0_value0 <= 0;
    layer0_value1 <= 0;
    a_buffer <= 0;

    layer1_value0 <= 0;
    layer1_value1 <= 0;
    layer1_value2 <= 0;

    layer2_value0 <= 0;
    end
    else if( i_aclken ) begin
        shift_buffer[0] <= shift;
        shift_pn_buffer[0] <= shift_pn;
        f1_ln_buffer[0] <= f1_ln;

        layer0_value0 <= layer0_value0_full[84:52];
        layer0_value1 <= a / 3;
        a_buffer <= a;

        layer1_value0 <= a_buffer - (layer0_value0 >>> 1);
        layer1_value1 <= layer1_value1_full[64:52];
        layer1_value2 <= layer1_value2_full[73:52];

        layer2_value0 <= layer1_value0 + layer1_value2 - (layer1_value1 >>> 2);
    
        for (i2 = 1; i2 < ITERATION_NUM; i2 = i2+1) begin
            shift_buffer[i2] <= shift_buffer[i2-1];
            shift_pn_buffer[i2] <= shift_pn_buffer[i2-1];
            f1_ln_buffer[i2] <= f1_ln_buffer[i2-1];
        end
    end
    else begin
        layer0_value0 <= layer0_value0;
        layer0_value1 <= layer0_value1;
        a_buffer <= a_buffer;

        layer1_value0 <= layer1_value0;
        layer1_value1 <= layer1_value1;
        layer1_value2 <= layer1_value2;

        layer2_value0 <= layer2_value0;
        for (i1 = 0; i1 < ITERATION_NUM; i1 = i1+1) begin
            shift_buffer[i1] <= shift_buffer[i1];
            shift_pn_buffer[i1] <= shift_pn_buffer[i1];
            f1_ln_buffer[i1] <= f1_ln_buffer[i1];
        end
    end

assign o_valid = in_valid_buffer[ITERATION_NUM-1];
assign ln_0 = layer2_value0 + f1_ln_buffer[ITERATION_NUM-1];
assign ln2_value = shift_buffer[ITERATION_NUM-1] * 55'd24973259072661437;
assign ln = shift_pn_buffer[ITERATION_NUM-1] == 0 ? (ln_0 <<< 3) + ln2_value : (ln_0 <<< 3) - ln2_value;
 
assign ln_value = !i_rst_n ? 64'hffff_ffff_ffff_ffff :
                    ln[63] ? (-(ln)) : ln;
 
//find the leading one 
assign index[5] = (|ln_value[63:32]);
assign tmp4 = index[5] ? ln_value[63:32] : ln_value[31:0];

assign index[4] = (|tmp4[31:16]);
assign tmp3 = index[4] ? tmp4[31:16] : tmp4[15:0];

assign index[3] = (|tmp3[15:8]);
assign tmp0 = index[3] ? tmp3[15:8] : tmp3[7:0];

assign index[2] = (|tmp0[7:4]);
assign tmp1 = index[2] ? tmp0[7:4] : tmp0[3:0];

assign index[1] = (|tmp1[3:2]);
assign tmp2 = index[1] ? tmp1[3:2] : tmp1[1:0];

assign index[0] = tmp2[1];

//calculate the sign bit of float result
assign ln_float0[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-1] = !i_rst_n ? 1'b1 : ln[63];
//calculate the exponential bits of float result
assign ln_float0[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] = !i_rst_n ? 11'b11111111111 : 11'd968 + index; //971 = 1023 - 52 - 3
//calculate the mantissa bits of float result
assign ln_value_shift = !i_rst_n ? 64'hffff_ffff_ffff_ffff : ln_value << (64 - index);
assign ln_float0[FLOAT_FRAC_WIDTH-2:0] = !i_rst_n ? 52'hfffffffffffff : ln_value_shift[63:12];

//adjust the output accorroding to the value of input 
assign o_ln_float = o_overflow ? {1'b0, {FLOAT_EXP_WIDTH{1'b1}}, {(FLOAT_FRAC_WIDTH-1){1'b0}}} :
                    o_invalid_op ? {1'b0, {FLOAT_EXP_WIDTH{1'b1}}, {(FLOAT_FRAC_WIDTH-1){1'b1}}} : ln_float0;

//judge if the input is valid
assign in_NaN = (i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] == 11'b11111111111)&&(i_data[FLOAT_FRAC_WIDTH-2:0] != 0) ? 1 : 0;
assign in_INF = (i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] == 11'b11111111111)&&(i_data[FLOAT_FRAC_WIDTH-2:0] == 0) ? 1 : 0;
assign o_invalid_op = invalid_op_buffer[ITERATION_NUM-1];
assign o_overflow = overflow_buffer[ITERATION_NUM-1];
assign o_underflow = underflow;

assign invalid_op = in_NaN || in_INF || i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-1] == 1;
assign overflow = in_INF;
assign underflow = ln_value == 0 ? 1 : 0;

//delay i_valid, invalid_op, overflow, to keep pace with output
integer i3;
always @(posedge i_clk or negedge i_rst_n)
    if(!i_rst_n) begin
        for (i3 = 0; i3 < ITERATION_NUM; i3 = i3+1) begin
            in_valid_buffer[i3] <= 0;
            invalid_op_buffer[i3] <= 0;
            overflow_buffer[i3] <= 0;
        end
    end
    else if (i_aclken) begin
        in_valid_buffer[0] <= i_valid;
        invalid_op_buffer[0] <= (i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] == 11'b11111111111) || (i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-1] == 1);
        overflow_buffer[0] <= (i_data[FLOAT_EXP_WIDTH+FLOAT_FRAC_WIDTH-2:FLOAT_FRAC_WIDTH-1] == 11'b11111111111);
        for (i3 = 1; i3 < ITERATION_NUM; i3 = i3+1) begin
            in_valid_buffer[i3] <= in_valid_buffer[i3-1];
            invalid_op_buffer[i3] <= invalid_op_buffer[i3-1];
            overflow_buffer[i3] <= overflow_buffer[i3-1];
        end
    end

endmodule