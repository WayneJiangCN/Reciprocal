//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
// Library:
// Filename: ipsxe_floating_point_a1_v1_0.v
// Function: This module is a lut for o_a1.
//
//////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ns

module ipsxe_floating_point_a1_v1_0 (
    input [8-1:0] i_x_hi8,
    output reg [51-1:0] o_a1
);

// o_a1 is the argument a1,
// which is in the taylor expression:
// a0 - a1 * (x - a) + a2 * (x - a)^2 - a3 * (x - a)^3 + a4 * (x - a)^4 - a5 * (x - a)^5 + a6 * (x - a)^6
always @(*) begin: blk_o_a1
    case(i_x_hi8)
8'd0:   o_a1 = 51'h59fb5ed31a53a; // a1
8'd1:   o_a1 = 51'h58f1113466024; // a1
8'd2:   o_a1 = 51'h57ebdb159c182; // a1
8'd3:   o_a1 = 51'h56eb99d60bebf; // a1
8'd4:   o_a1 = 51'h55f02c01834ab; // a1
8'd5:   o_a1 = 51'h54f97143f32f8; // a1
8'd6:   o_a1 = 51'h54074a5dad118; // a1
8'd7:   o_a1 = 51'h5319991830593; // a1
8'd8:   o_a1 = 51'h5230403b80169; // a1
8'd9:   o_a1 = 51'h514b2383f98ba; // a1
8'd10:  o_a1 = 51'h506a2798a4955; // a1
8'd11:  o_a1 = 51'h4f8d3201f7684; // a1
8'd12:  o_a1 = 51'h4eb42921077ca; // a1
8'd13:  o_a1 = 51'h4ddef42721e16; // a1
8'd14:  o_a1 = 51'h4d0d7b0dc5894; // a1
8'd15:  o_a1 = 51'h4c3fa68efa737; // a1
8'd16:  o_a1 = 51'h4b75601e00e22; // a1
8'd17:  o_a1 = 51'h4aae91e054151; // a1
8'd18:  o_a1 = 51'h49eb26a6fc452; // a1
8'd19:  o_a1 = 51'h492b09e82bd9c; // a1
8'd20:  o_a1 = 51'h486e27b9240e0; // a1
8'd21:  o_a1 = 51'h47b46cc85d714; // a1
8'd22:  o_a1 = 51'h46fdc657f0e2d; // a1
8'd23:  o_a1 = 51'h464a22383dd97; // a1
8'd24:  o_a1 = 51'h45996ec2caf3b; // a1
8'd25:  o_a1 = 51'h44eb9ad55df94; // a1
8'd26:  o_a1 = 51'h444095cd489dd; // a1
8'd27:  o_a1 = 51'h43984f82e77ad; // a1
8'd28:  o_a1 = 51'h42f2b84550d97; // a1
8'd29:  o_a1 = 51'h424fc0d63105d; // a1
8'd30:  o_a1 = 51'h41af5a65d2067; // a1
8'd31:  o_a1 = 51'h4111768f4cac8; // a1
8'd32:  o_a1 = 51'h40760754e110d; // a1
8'd33:  o_a1 = 51'h3fdcff1c74a83; // a1
8'd34:  o_a1 = 51'h3f4650ac34349; // a1
8'd35:  o_a1 = 51'h3eb1ef2757ede; // a1
8'd36:  o_a1 = 51'h3e1fce0b08548; // a1
8'd37:  o_a1 = 51'h3d8fe12b62323; // a1
8'd38:  o_a1 = 51'h3d021cb098630; // a1
8'd39:  o_a1 = 51'h3c76751432116; // a1
8'd40:  o_a1 = 51'h3becdf1e64213; // a1
8'd41:  o_a1 = 51'h3b654fe38496f; // a1
8'd42:  o_a1 = 51'h3adfbcc196d64; // a1
8'd43:  o_a1 = 51'h3a5c1b5defa2c; // a1
8'd44:  o_a1 = 51'h39da61a2efda4; // a1
8'd45:  o_a1 = 51'h395a85bdd4ee7; // a1
8'd46:  o_a1 = 51'h38dc7e1c9e2db; // a1
8'd47:  o_a1 = 51'h3860416c05f8e; // a1
8'd48:  o_a1 = 51'h37e5c6958e0ce; // a1
8'd49:  o_a1 = 51'h376d04bd9e12a; // a1
8'd50:  o_a1 = 51'h36f5f341b3b00; // a1
8'd51:  o_a1 = 51'h368089b6a3608; // a1
8'd52:  o_a1 = 51'h360cbfe6e9616; // a1
8'd53:  o_a1 = 51'h359a8dd10a091; // a1
8'd54:  o_a1 = 51'h3529eba600e78; // a1
8'd55:  o_a1 = 51'h34bad1c7be139; // a1
8'd56:  o_a1 = 51'h344d38c7b114d; // a1
8'd57:  o_a1 = 51'h33e1196560da3; // a1
8'd58:  o_a1 = 51'h33766c8d10396; // a1
8'd59:  o_a1 = 51'h330d2b566e75e; // a1
8'd60:  o_a1 = 51'h32a54f0353558; // a1
8'd61:  o_a1 = 51'h323ed0fe864d4; // a1
8'd62:  o_a1 = 51'h31d9aada9057a; // a1
8'd63:  o_a1 = 51'h3175d65098086; // a1
8'd64:  o_a1 = 51'h31134d3f4778e; // a1
8'd65:  o_a1 = 51'h30b209a9bbaaf; // a1
8'd66:  o_a1 = 51'h305205b67d04d; // a1
8'd67:  o_a1 = 51'h2ff33bae808d5; // a1
8'd68:  o_a1 = 51'h2f95a5fc31928; // a1
8'd69:  o_a1 = 51'h2f393f2a83697; // a1
8'd70:  o_a1 = 51'h2ede01e40af88; // a1
8'd71:  o_a1 = 51'h2e83e8f21fc16; // a1
8'd72:  o_a1 = 51'h2e2aef3c0423c; // a1
8'd73:  o_a1 = 51'h2dd30fc614928; // a1
8'd74:  o_a1 = 51'h2d7c45b0fd7b2; // a1
8'd75:  o_a1 = 51'h2d268c38f79f4; // a1
8'd76:  o_a1 = 51'h2cd1deb50aa4b; // a1
8'd77:  o_a1 = 51'h2c7e389655a0d; // a1
8'd78:  o_a1 = 51'h2c2b95675d692; // a1
8'd79:  o_a1 = 51'h2bd9f0cb60729; // a1
8'd80:  o_a1 = 51'h2b89467db00d3; // a1
8'd81:  o_a1 = 51'h2b3992510eca9; // a1
8'd82:  o_a1 = 51'h2aead02f13e03; // a1
8'd83:  o_a1 = 51'h2a9cfc179358f; // a1
8'd84:  o_a1 = 51'h2a5012200ae92; // a1
8'd85:  o_a1 = 51'h2a040e73133d2; // a1
8'd86:  o_a1 = 51'h29b8ed4fd5991; // a1
8'd87:  o_a1 = 51'h296eab0985a3d; // a1
8'd88:  o_a1 = 51'h29254406df388; // a1
8'd89:  o_a1 = 51'h28dcb4c1a81ab; // a1
8'd90:  o_a1 = 51'h2894f9c6356b6; // a1
8'd91:  o_a1 = 51'h284e0fb2f4bdc; // a1
8'd92:  o_a1 = 51'h2807f337f8ac6; // a1
8'd93:  o_a1 = 51'h27c2a11688d0a; // a1
8'd94:  o_a1 = 51'h277e1620b4fef; // a1
8'd95:  o_a1 = 51'h273a4f38ebabd; // a1
8'd96:  o_a1 = 51'h26f74951935eb; // a1
8'd97:  o_a1 = 51'h26b5016ca7194; // a1
8'd98:  o_a1 = 51'h2673749b55988; // a1
8'd99:  o_a1 = 51'h26329ffda35a0; // a1
8'd100: o_a1 = 51'h25f280c20f4bd; // a1
8'd101: o_a1 = 51'h25b314253a11e; // a1
8'd102: o_a1 = 51'h257457718fcbe; // a1
8'd103: o_a1 = 51'h253647fef4457; // a1
8'd104: o_a1 = 51'h24f8e332717e0; // a1
8'd105: o_a1 = 51'h24bc267de8747; // a1
8'd106: o_a1 = 51'h24800f5fc4242; // a1
8'd107: o_a1 = 51'h24449b62aea1e; // a1
8'd108: o_a1 = 51'h2409c81d4846a; // a1
8'd109: o_a1 = 51'h23cf9331e0d86; // a1
8'd110: o_a1 = 51'h2395fa4e32a0b; // a1
8'd111: o_a1 = 51'h235cfb2b1f619; // a1
8'd112: o_a1 = 51'h2324938c6f196; // a1
8'd113: o_a1 = 51'h22ecc14090884; // a1
8'd114: o_a1 = 51'h22b582205b686; // a1
8'd115: o_a1 = 51'h227ed40ed44bf; // a1
8'd116: o_a1 = 51'h2248b4f8f2145; // a1
8'd117: o_a1 = 51'h221322d564f4e; // a1
8'd118: o_a1 = 51'h21de1ba45ef70; // a1
8'd119: o_a1 = 51'h21a99d6f5df1e; // a1
8'd120: o_a1 = 51'h2175a648f6ec7; // a1
8'd121: o_a1 = 51'h2142344ca2dd9; // a1
8'd122: o_a1 = 51'h210f459e8cc03; // a1
8'd123: o_a1 = 51'h20dcd86b60f1e; // a1
8'd124: o_a1 = 51'h20aaeae81dd0f; // a1
8'd125: o_a1 = 51'h20797b51e591f; // a1
8'd126: o_a1 = 51'h204887edd1420; // a1
8'd127: o_a1 = 51'h20180f08c4eeb; // a1
8'd128: o_a1 = 51'h7f40eee939a6f; // a1
8'd129: o_a1 = 51'h7dc852da66383; // a1
8'd130: o_a1 = 51'h7c56ea38dcece; // a1
8'd131: o_a1 = 51'h7aec840c0d24f; // a1
8'd132: o_a1 = 51'h7988f1045cb2a; // a1
8'd133: o_a1 = 51'h782c0369ae4bd; // a1
8'd134: o_a1 = 51'h76d58f0abfc5c; // a1
8'd135: o_a1 = 51'h7585692d542eb; // a1
8'd136: o_a1 = 51'h743b687f1e972; // a1
8'd137: o_a1 = 51'h72f76507630d6; // a1
8'd138: o_a1 = 51'h71b9381943f20; // a1
8'd139: o_a1 = 51'h7080bc46b265b; // a1
8'd140: o_a1 = 51'h6f4dcd53f91ec; // a1
8'd141: o_a1 = 51'h6e20482bd97c6; // a1
8'd142: o_a1 = 51'h6cf80ad433278; // a1
8'd143: o_a1 = 51'h6bd4f4632f073; // a1
8'd144: o_a1 = 51'h6ab6e4f4e6ba7; // a1
8'd145: o_a1 = 51'h699dbda1822fc; // a1
8'd146: o_a1 = 51'h68896073c54ff; // a1
8'd147: o_a1 = 51'h6779b060080ce; // a1
8'd148: o_a1 = 51'h666e913b93766; // a1
8'd149: o_a1 = 51'h6567e7b45ec66; // a1
8'd150: o_a1 = 51'h64659949279d4; // a1
8'd151: o_a1 = 51'h63678c41e0ee3; // a1
8'd152: o_a1 = 51'h626da7a874585; // a1
8'd153: o_a1 = 51'h6177d341d1e83; // a1
8'd154: o_a1 = 51'h6085f7874a750; // a1
8'd155: o_a1 = 51'h5f97fda03100e; // a1
8'd156: o_a1 = 51'h5eadcf5bbfb78; // a1
8'd157: o_a1 = 51'h5dc7572b3d53a; // a1
8'd158: o_a1 = 51'h5ce4801c5fe03; // a1
8'd159: o_a1 = 51'h5c0535d3e9f4a; // a1
8'd160: o_a1 = 51'h5b2964887fb08; // a1
8'd161: o_a1 = 51'h5a50f8fdb0e21; // a1
8'd162: o_a1 = 51'h597be07f35e3c; // a1
8'd163: o_a1 = 51'h58aa08dc5cde3; // a1
8'd164: o_a1 = 51'h57db6063a53aa; // a1
8'd165: o_a1 = 51'h570fd5de872ef; // a1
8'd166: o_a1 = 51'h5647588d65678; // a1
8'd167: o_a1 = 51'h5581d823a6ec9; // a1
8'd168: o_a1 = 51'h54bf44c3f7799; // a1
8'd169: o_a1 = 51'h53ff8efcac939; // a1
8'd170: o_a1 = 51'h5342a7c44dc1f; // a1
8'd171: o_a1 = 51'h528880763e5f7; // a1
8'd172: o_a1 = 51'h51d10acf878fb; // a1
8'd173: o_a1 = 51'h511c38ebc0f54; // a1
8'd174: o_a1 = 51'h5069fd4216d5e; // a1
8'd175: o_a1 = 51'h4fba4aa26c6c7; // a1
8'd176: o_a1 = 51'h4f0d14329935d; // a1
8'd177: o_a1 = 51'h4e624d6bc0158; // a1
8'd178: o_a1 = 51'h4db9ea17bf3c2; // a1
8'd179: o_a1 = 51'h4d13de4eb7c7f; // a1
8'd180: o_a1 = 51'h4c701e74ac228; // a1
8'd181: o_a1 = 51'h4bce9f37342c5; // a1
8'd182: o_a1 = 51'h4b2f558b46505; // a1
8'd183: o_a1 = 51'h4a9236ab14a57; // a1
8'd184: o_a1 = 51'h49f73813fd4dd; // a1
8'd185: o_a1 = 51'h495e4f848d4c3; // a1
8'd186: o_a1 = 51'h48c772fa95128; // a1
8'd187: o_a1 = 51'h483298b14e13d; // a1
8'd188: o_a1 = 51'h479fb71f90ace; // a1
8'd189: o_a1 = 51'h470ec4f619bd7; // a1
8'd190: o_a1 = 51'h467fb91ddf558; // a1
8'd191: o_a1 = 51'h45f28ab673de3; // a1
8'd192: o_a1 = 51'h45673114772ee; // a1
8'd193: o_a1 = 51'h44dda3c01504a; // a1
8'd194: o_a1 = 51'h4455da739056f; // a1
8'd195: o_a1 = 51'h43cfcd19db0d6; // a1
8'd196: o_a1 = 51'h434b73cd399b6; // a1
8'd197: o_a1 = 51'h42c8c6d5f2108; // a1
8'd198: o_a1 = 51'h4247bea9062cb; // a1
8'd199: o_a1 = 51'h41c853e6f8106; // a1
8'd200: o_a1 = 51'h414a7f5a9921b; // a1
8'd201: o_a1 = 51'h40ce39f7e2c66; // a1
8'd202: o_a1 = 51'h40537cdad8949; // a1
8'd203: o_a1 = 51'h3fda414673a26; // a1
8'd204: o_a1 = 51'h3f6280a3969dc; // a1
8'd205: o_a1 = 51'h3eec34800a5ae; // a1
8'd206: o_a1 = 51'h3e77568d828ad; // a1
8'd207: o_a1 = 51'h3e03e0a0aa4f3; // a1
8'd208: o_a1 = 51'h3d91ccb038619; // a1
8'd209: o_a1 = 51'h3d2114d40a8a2; // a1
8'd210: o_a1 = 51'h3cb1b34448235; // a1
8'd211: o_a1 = 51'h3c43a2588b68f; // a1
8'd212: o_a1 = 51'h3bd6dc8711575; // a1
8'd213: o_a1 = 51'h3b6b5c63efde3; // a1
8'd214: o_a1 = 51'h3b011ca0522f8; // a1
8'd215: o_a1 = 51'h3a981809baf35; // a1
8'd216: o_a1 = 51'h3a3049894c2d0; // a1
8'd217: o_a1 = 51'h39c9ac23149f0; // a1
8'd218: o_a1 = 51'h39643af5627da; // a1
8'd219: o_a1 = 51'h38fff1381b41d; // a1
8'd220: o_a1 = 51'h389cca3c186fb; // a1
8'd221: o_a1 = 51'h383ac16a8925f; // a1
8'd222: o_a1 = 51'h37d9d244584cf; // a1
8'd223: o_a1 = 51'h3779f861973d8; // a1
8'd224: o_a1 = 51'h371b2f70ecb96; // a1
8'd225: o_a1 = 51'h36bd733708112; // a1
8'd226: o_a1 = 51'h3660bf8e18531; // a1
8'd227: o_a1 = 51'h3605106547628; // a1
8'd228: o_a1 = 51'h35aa61c038d51; // a1
8'd229: o_a1 = 51'h3550afb68c77a; // a1
8'd230: o_a1 = 51'h34f7f673645ca; // a1
8'd231: o_a1 = 51'h34a03234ee54d; // a1
8'd232: o_a1 = 51'h34495f4bf0b86; // a1
8'd233: o_a1 = 51'h33f37a1b5a641; // a1
8'd234: o_a1 = 51'h339e7f17d5cfb; // a1
8'd235: o_a1 = 51'h334a6ac75f262; // a1
8'd236: o_a1 = 51'h32f739c0dd451; // a1
8'd237: o_a1 = 51'h32a4e8abbd8e5; // a1
8'd238: o_a1 = 51'h3253743f92729; // a1
8'd239: o_a1 = 51'h3202d943b4a13; // a1
8'd240: o_a1 = 51'h31b3148ee6c6f; // a1
8'd241: o_a1 = 51'h31642306fbc80; // a1
8'd242: o_a1 = 51'h311601a07f611; // a1
8'd243: o_a1 = 51'h30c8ad5e611d6; // a1
8'd244: o_a1 = 51'h307c2351a18e0; // a1
8'd245: o_a1 = 51'h3030609901b2e; // a1
8'd246: o_a1 = 51'h2fe56260b4823; // a1
8'd247: o_a1 = 51'h2f9b25e2127f8; // a1
8'd248: o_a1 = 51'h2f51a8634f51d; // a1
8'd249: o_a1 = 51'h2f08e73731495; // a1
8'd250: o_a1 = 51'h2ec0dfbccac61; // a1
8'd251: o_a1 = 51'h2e798f5f3571e; // a1
8'd252: o_a1 = 51'h2e32f3954f3df; // a1
8'd253: o_a1 = 51'h2ded09e17918e; // a1
8'd254: o_a1 = 51'h2da7cfd1574eb; // a1
default:o_a1 = 51'h2d6342fd9386f; // a1
    endcase
end

endmodule